��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛������^���P�C����L�9jc��?3�8*���	̆����=H���Wݝ�QE���o��d)J�%����e���vid��:�x�y��d|W̱p�)^�MJ��Ǟ�H� �a�C�����c�&�|�ۣ"�6����=a�BT7�](���~�՜�l�ܞ&�f:XΕ�B�:�,=��Q9{Våi��}Q(:&o`�G�5�e^�5���3�n���� �c��1!Hz�'�<~23�wt�u)J��[�zN-ю��4���)K|F%FGU�� UwՁ�^������b��t ���*�$|����]w8�M�:�02����/n����X���<LY�|���_n��i�DlҬG�	�P��,��܍�����Q��m=_������뉆BNO9Zh&�Z �S}.v�������Y�UL���i�F=|�7��E5��\��o�q�L[/*LG6D!u4X^��H�8装it����M�	�[�Q��E$u�ht"!?�"ab8��Z�2{��=0��F��o(K�2��|���	y��DVM����t)�xC;-���AI��_���bމy���y��B��c�6j��y�빌��K�Lo������@Odt�`0W<�-�ۊɹ���$X���?�q��o\3��GK
�3?�v�Z����B�ǧ�\�q]��e��f����p�e�}��ג=�9&�;�E�ǋK�L�lE��E�>���X��'��i�
4w�!���f]������us= -D8����&�x�3J�8�v=�jI,j��_4�խ8��?ߕ�);�Fզ�=ժfu1�u�Q0��Y���;+H8t�<R��Pc�/��NsإG���K�Ê�<�%��X 5S�O�bEdL�)�'���OR�MW�uK�I�E��/e��>Y���0s>(��*�]�zX
�f5�&����a�?���"����Y�U�u	$����ް`'as��U��5H�\4�0㭛��4�?6*��d>N=��_�2�M�D�l�U�20�	"��2��aP{��k���i����w��M�)��:+8=�N�+�.;�|�f-ߎ���*lSˁB�^~x5%����F�������b1%��[��c���	}h�<���m�~��#g��T��Y=�8\�[/�t��\`�<l����@���^�9��~z(����F��j e�规�V���ܬ��j�졹*��,պ�(�ߴ����C����L�G#��
G@nm�����|�x���S�۵�%~��ü6	j�	��2�I,��}�S�Sp�H�\if؉���˻������zq
1�Pk��,N繙=ߒ���<!O�y����O��E.�.�ry�y�?���d�>�2��P�-�ߎ�q������o<���5��?-/��iw�B��w�:&���O9��K��� e�@��0��&�ݰ�b���(eG�Al����\�,�,��F�ЪfW9�6S��#�%�:Vu,ա�5�����[�[�=�3�5���������٢v�j8p���*�$ܠ�Ӻ����4�2N;?�u�My��7p| \���[�w�*�ơT�ċ�����F��\��̀TS�D�G_����L6�R��H/k��P�{~��S�B�sՁ�T�|`~.�/��&�B����S]������I���f~I4����� �s%�����m�N�v]l��eBaaȤJ�|>I��N��Q�)���-Ǩc��`��R�������XO��?��}>+ʑ��������r�ƿ"�R�K��5*"�i��z��s��9@1Vv�4U��E���g�Z.�n������b:M"k_K��[�s�q&0��;dK��a�X�����q��eZT�:m���6�T��T�ڙ*!Զ�����9�1uZK!��)����&\�f�;��=�wZÉ7)�Q};LH3�߻n�c>�������j�a��"S^U��³����|��Ō�t��h��ȀY3�0��t�w��.�!���z-	��gr��3�[�� ��'���%�5���[i	���Kuh�X^y=�@	���/�xaXc����7l4���Hett��>v	��vCc�(4R�c�bA��27��&+l/JY�	��h�s�8"	J���o<�<�h�Ո����A�I)�b0���t
k�'���M~n��0S���M|��5�4i`/3��	�EΑ���@�DʉIDf�O̜�䞶3jc�����>"�|z\�G�>��M%�7ěbF�_a���*H�-_�;2��ǚ���#��[�2�.3�m�m��d79���k���� A��VM�|/5�%�@�5kK2m���V�P5�_8�S���h�-'���"�N�m=0{�Tc">�4�}���8��+�{�E��`p�A�����+F�'��f�.>E;�Q�*���(��H��xFz��)��듡�=�>�󕣁˼� kY	�v�?߼e�e5����\UJQ�(&��. �✞�%]":�ý�u�:k��	Ώ�h ��W�DM�mмj������l���%��"���0�uXJ�H���-��Hf��@�N�a/���V��-8���Ę����?�p�I卉mq�u�`�񮿱(�o�;	��SAt�%��4N���~֗���f����CS��V0*I�����k ��:�V�o�� ^�`E�HkbnX�ˢS����2o1ޛ����Ū0L��t[��[{�x�Ľ1b�$>�yq)�X¿'+�����Ъa� ]�R}x?��{�qW� ('R��U�mU���$#���\�(k���I"Xu'SC�.��ٵ��_c�+��2������e�H�����)�r[X�f�oTx�����0�'��9Gm�yǑh�Ԉ�~Q�fo�_a��f�dIV����m=M�3�Wާ����;�W��g�]�Є�u�
e4�rPz�y����K�}���y�jI�_o�.�fQ�ր_��g  �2�d#j�B��j�ny�����q�=K����Z�Cd�T��Uq=:0B��xM��)�H�(y;b{e�����<1��^Ɓ�
j?Gr��e$Os�98����4J�(����׬p��9:���7�A�,����]d<6	'��a���A��:��{�r�GCu��~Lʰ���T�\4�dɁL�����r��H�	��ؗ�xX�����DLuZ�:�W(� ��
IbZD��� ����#të��J��}
��\D`�W�Ҏ�Z��05�#e�/�A�yv&��r�*ٞ�hO���{��b�$���ǲ�	��~�����(�	rF��XxcT%R�黹��>oS���lX���`=g8*F�y)�]��!xL{��Xc���>�ς	������kLn�Q�nJ���-^�"���+�<$����Q�)��f�aW9��2_rp��4akJeS��3��Um_��sv/��o�)��ʽ<Y���f��4��	Xo�Oi�;Xf��piʟLY<
Q_lNL�P�W�YN�;�皽�'@)�����w]&~A2�o	&u���%�5*6jlyɱ8��x:�f�=�=S��
�]�*A�@2L���A�[�����;^��7j;(%b�S��c��3�]�S0�g��/��P�3G6�M��s��T��r����$Cۋ�`'@�i�M�[P�P�s�]��)ZP�s��T@��8*��ٲ!�ﷸϠ�F��5<��B]����꩚-���jl�z��I�	�BƯJ@�ȝ~j�5`w��9�/]��-���\w����cO�S$Ψ21����CN��4o��T���*�|�Z�,(#-g5B��3����7��(u�]ITj��;�&�c�̄x$����
�ۤz��L���a��4�[�@~�3��!�D���n%%J��@S�4�_��q����n�GN�����#D�1��\����V��]���>D��R����9Ov~0��]�LwY������<��x[�jA�RMZH��-k��|z�'(7��y��,e>�=��:���n�%�:�:���)+�Zy���~��l=Zb���K��DD�@=��E���ȼI �rж�ྲྀv'~��	���,�8}���ܩbc���Ng;]�Y�����Fr�d�X`�ʄ���2j�z�H[���&S�P�2k�lT
���x[Jj�<�����4@}e���ZR�}z����orH��%������p�uK&ͨg3ں_�{s���4 �T��2�ͼ{I��6���7b��&Ď�]-4~��~7�_�'�|N�\\ Z�ý����lqg#��e�����rP<��A���w_(�K�G����S+�hg��ќ5��\�.~q�%��I:Ydm��Dz��V����Nm3z����_[�ܾa�	�!B"�4���*�[O��V�j�Uu������I���凰��y�)m88��LZ{�<�F�<WGF4���!�"��;���Ds��"B���j���}�ɠ���W�C��PR！f%)
�:���?��R0G��`3�OI��b��� Bc��[��r�b�bʂ�� kK��ˉ�ڴRƖ�DX����(�9�o�y�]�W\}]�uo�I_?u�$у�q@{4�^��g'�4�.�D;���џz~�>B���	Q��!�Q/�}��>�Z ����uS�g�\�b:�Ǯz�FP��q^��`�cf��\�Uv�*/0<�nt�(�E�|N�`��h��ٷR��Q�p���O��gJ�E�}j��ð	3�ȿX\��}��_�1���P�F��R��6��q-y��Z� ��{�#w7�Kz������d:�_��Yg\zL��������v����.詰7۬���\�B;��ae���}�P��φ�X�Ф�\�^6�_�Ii8p�ҽ�L�>��Jr�6��D{�,�:Q�?a0���6�n��t��3�j�%g�C�Gr��-쵆�;��eQ0�����Up�)��&2x��Z}t��\���Ps��B>��I�Ӯ!w�]��R��~��N���Vyv��ߘ'�y��5	O���p�T5؝l0�s8ʔ����:�x#SpY{�������~M�s'�:�Q }Ӈ~:�%�g������
� ��6�<�+��s�N������-m�i�D�b}���}��w;�؟9{̚�E�i˾���9fZ��á��rY{��	W=aiV��.H�̕#�$ѾW[)�mt���BH�� �E�X�a��z$�wY Ok�2s,�>�h{�U{����n�e�?����t }�P�s~_��F���Б�J��lH�Y`����-��mF�����ş�������"G���K�Q4&~i�{�ej%���K�C��b������v�b�-�QY���B�p�X�{�eE'T�t���ɣYO���Q����@C�}���մ̆�li��v���>÷4:��*l{�ȟ|ң�ESWG2�5��j�Uƃ�ѓ�)�~�!�'��o����βV�ܸ�j9h�pF�Ow}^l�,?�b�~x�t�<������37:y��>д/��@ں�87c?�x_�l,���� )8��=�̖�v%�A�s)O���'B8S�Jp�k��D^k;�Gga�<�E�	o���C_2l��F�?Ӳ�9~1 1����ˣ�FC�ke¿ʜ�8(��n}���"oB�,�~�vi�	\����������f���wR�і�x�S�������+�}�Q A�y���u��
cw��='�/.�/>��� �&S��5�*�ti�P��Eu�!n��)E��H�<ԁ��L�ŵ)��T_��ݒ�mU�k����<����G[>�X�i#��h`s�=K}rS� �@���Wz��r��rP�(���oP�==��݀8�ʹ��w��g>s֓�"�����d`7��%�u����h��d4C�[1���q�ʎ'[N|�n���U��IR�c��Oc+XNn5&�K�Cnw������A�jG�)����Y<K�zޔ(�<�a���\ou��1$��t�������}�)�"	�#ye=�
�E\[���)�x'Hj�Y��c�); �	Uv����"'��=G;�ͦm
,�X�fQ�h343�����������A�wI��z3U:���婯'n)��壘�?$ ��
������X(���̄t��w���!��<7�� �Ί�xj���� �)(J�Iv���bd���N��g��1	>�_ ���XK�
 ���?�^��mj���0ĸRgH�c�0�#�D}r�,�-�A�x���3��,���H���FC!�oY����{b��!$����И���Z�&��FD�-ȍ�[�s���� �6�W	~���?�֯�ܐП�	V�ꄉC���x�!/���o��ݏg�Gf���v��GT��3�Bc��2����K��3� _�e�U%�R�g�Ⲽ�y�&ۀ��kh�M���|���;����������MI)�rJ�����\������+�I&��	���֘��۫���0k$�����;/���}��0Y����5܅ˈ���W�X)+ьR��Pg����w}=��;ח+M������@��߮��,�Xa5�k�o�V}���17?��'�(�yWbjeԐ^v����G�4�8�LIhPx��-ۥ������D�>�����]?a�𪧈����)��p��z�>:Zhɋ��	t��~��fO:,_���|R}x�*pvw����/�i4t��@����$Z�H�rI�d�(�n3��HƘ�8����̯ �����G�xp��\uX�i�'B-lR�)Q�C��S�"��Cb2Ae3�h�YV�#��?� J��(ޯUe��ge,�E��A	T:I��1��~ �`����t���7�E��_�w���d2��qZ�r��$d4��&ckZ�R,�r�e9�nMi��� �]h�^M��$Lh4���a��2�Ï��G��	����9oR����z��wşA�ǀ9�t��i��& �\X,*a)z� �fQ������!u+
��A�95p�fL���dD�lVw�|��q<������\6�U��p���[�qY����sg��^2Y��j�(5k���"��s�P����y��닼��.�MC�h�Z�T�C���빻j��MnT�o$?��.�^~e$y�O�F�S��_�ܑ���A��3j�N�TI����Ѓ�����K��D�ny����|n��k+>q��W�� |�z��{�K��^�$��𰴽�0�)�+��8k�XN�Z"^��'�'���=�6��;��)4r���K�{J����F�j"��vv>���~Y(n�
Aځ��Qn��i�7��x��{�7U��Ӻ�uGDA����B$A9��:���!~�Qk>=3Kط�a�7��[��8a5N�T7�U�©����8��h�%R��N�ZC�"f��_��r� E��.�S�# *�RA��q�Q��k�0��,�/��I����ٺF[��������_6B16c���9*Ղ
�|Cn$~�V��Ą9f�ݻ�,����Էp{ ��L���*������SG�G�]n[��XV.c<�� �(O��C��}��� �P�p��!�g����y�$ɂ	N���C���l�펯|C��3E���`!A���^5\�^�A�כ0hZY~����uL�p$��ޝ����=k�KD.�t+�?��} �0
G{�ET	��+��y�o��^�>� 5�bX_�ң���P�9y"���*��#���h���Ş4����YN|�X�Ur]��m����uM�!�y(A6݆#�xcD��x���2�(�/w���������$y�г��g6���ݳp �K/!���n��r\�F���Ǜ��hS}м�R��5���L�6��{ެ}[9����$�1~�Эqz�R�(�p-7�?�N���Q)3��g�dY13�&��W9_UT�_�Cz c�b������U09�ͥ~w��r+��,J.���H��ί�F��jf�HNT���?��
��.�u�1*�w��۸��s�i���Y�ɑ�����w���Qn��d�{�-���|n?�Ԑ����FDgk����je?ԋ8�5�-����vC����u�;�~4C=�D�?S���~�6V�>%��=Gf�)#*��:Roam����ytF���+���>� R����������Rz5��������}7�U��wj·�G��R�s�Z��!$�������g����〢�H�'�D�����䖱΁W�j_ڭT��G!�~Y�qDS�������s�px_�g�8GL����q��f�$=К�s�<�f&�-��'��o;�������k��C�� �ȸ ��Y�C7o�:#�s��Y��iX���&O�'!�ݡ�7ڀ!C"P,�=�eh0��>e��c'ei\��
��H�r�{�%�r������>f(ϣ���m@����;#W���*5Bc�H}��X�& A%����(�3V.���QO�MB���:�в���<��[�B�'y ֓v}�wb؈0�h+ĉ�, cY����٠d�nC�������Q����hn��x���,e�e�7v��~�
M>w|����x~tI�ZG=�����N,��#z=���k����!v��`&A��F7�p��Q�x3�t� y�tl$�,"�ZF����'���J�|]{�@xs��M�'5�Bj����WemJ~�Tb��P92j�jۉ!���
k�ݨCo6�S��"xB��Y;�eLCD)!��ġ�C�ʸ:d�{p���]8.���h�P�dPs�.�o���aa�oMZǣ3�6���3�Vyd�L��7Xi��7��G	%���+���r.���ώv�����΃�:���%s!�%�ezɤFVl�:�fR��eYT�;Ѻ��uV�m�a W`(��mgMk����\Mv���wd։z�'�c�u�vKQ�HR��)mX��j���9��w�`~�;��]Jv��8�=h�z�5+#��؀�� 6nM�8�4�O��n���߸}�aG��P�"C�`z ��RW�Ճ/�弳����܃A�qS�Dq>�)���pq�5o�*ܥ����քo#�f��wz�����90w��A(;��]$w��%�=�jI�E76*RsB���C!flѶ�^�|TYI�I�<��h�g}��}/0���O�G�5{���?o��$Ep��Ʌ�@~pҸ�'g�as��&�o!��� $�:Q?����`\���W���@���@��~E	���T�'q���C����;�PiR`>nK�,�	��)�����ͯ|C rRR-���L]۩�����0H|�h�|�z~��Ld ���
;@�fZ9�/��z6��˺x����Z�� C����cQ �4�9�������8���yAb`�M��5�n���J����~�s��3c<Q��[Ȑ��i���r����]-e#��ks��4�w���x���I����)�e�f�e��i^J��u_��+������4�*`���\d��C�@?�c���/\�2'B�,����:97S3V����PH��򓵎\9�X�.�m{/>m2��$���P��@�a
�U7�N����^�R��B/�y���Ң)�%�}I���D% �?��u��=�c�czW�����@��5���|R%j������?J�S����t�L�`oT��#����^(��P�����tlu�4Ft�hƈ��0�7�0���aV6=�x��ەQ���ڠa��J�+��I;���-rQ4�x'R��(Mp��DlG,h�I�"~a�V�򽰀[���H�9�l�}�=���I����� [T`����9$�Vֱ�-:�����Y�h&G�(zs�FG�(�)��M'j��ױl�Y���Z�{��ㆺ��F�2X�B��[�� (��Y��:�ifjC �=���q�@>����B����9�[�q��Ů�=w0᳣_T�B>*k����y��sܔٳ�M��gk�nlW3VY��e�z.����O|�śQԼz��|v�����<"�Ц��	P��:f,�c�2!�>�]���t�9X/��/8�3v�Z���i�_�+�^d��6��u;���bگ��୸s�a&d��d�0��v�� (\C�G_�y-�}�l
���7&�@5ܭn҄i��較��d���e�[���R�a����x��߉:c��oP�����C*�M �D-��n��CC4~�p ���?� �[%�%�1+���ʝ��g�?�
.VL�K����ڱ���!RȲ/��~�YJ��x��������h��᰻��ܰ\)�F�u$ ^� �D&���`�X�j(�+����K����6�����������w/�"65X����QΈ��!�
�&Qg{��1��ޱ�����G?�������k������%��a~aUF�f`�o>�(��cECa����[y���d	oU+��N)!y�2P?�[�p��?{�-�{"��o�#��#�'��
��P��W4f�o��q%c)P�ì@^�Ue��}V�����M����H��yʿ���r(�f9{0ܑ8�s7��j
KM�	a>
�H�?Z\.Z�_�u�N�Ċ�r`�t*}���BRd�y�i@4"���},{�Xoq�7 �lĞȺ��g#􎒸� ����ח��b��>M�ܾ�.��]GM4�mf[���5;�!嗵�\nU]�����ߪR��ɘ��2��N���(� �q���E`��f4s"�����k�v�������)L���%���rlx�9O'�F �H+)@p�u،�f��a\+��d����qa�B����m��Y��6�>����Q'HM7����)�?���F�MT4��/�*im���'�$vsib��=�/�I��"[��7*�r�j���;��h�d�ҭ���;�Bt
P�<���r2������0�a���EbX]�������]^��M��2/�C�mUe��*6!>�,�	n�a���X�/:���e+��fJ`���g�R$��+�6�x�b�|��[Mƀ��ϡ���B�[BAau.}�9���%��l%���0���(pr+kw[H���}�����hW�O���ṑ;�).Cױ:d�>#PW53���:%c�Jk���C㽹��H�=��I �S������~�V�
����Щ��+q���m�)�kOw�C5Ē��sF���nhնR��ӗ�[�ӄ<�F��E��-ݿXFz*X��{	�ι� k��TI���ܱN�vH�8ۼ�:X��-Ӊ=� �JЮ>Q��)�z?� Eb��:6���B'�Ý��q]�A�+��Q�������0{z��7*!��4����AbwCr�x��Uy�GK����k'`֢�K-�N����wx��ʫ�'�< t�e	͸QB�\�8Hc�tи�0�n)vl��1�	@�@r���I 7�θ�De6
g8W���9��C{J���=a������^���K{��Yq�F9��A�VQ�0Oy>p"����G]�w.����")t둏ѱ5���/���W%p���mH4��+|O!�܋W0ʓ>�������U��~T��5Mg�� �ݻ�g;�ٗwuk��7;���	����µ?��xz.SRt��"�f|������"z�}��0�	�����Z����Y�J�V��8�uvp~��Ws;B�����g�z)��-�ͨ׫$�:���F�;�z��Em��3��H�dh��A�`����p���ݐ��?_Fx�IM��O�����S�|����?!�X�z��S�u�o��l�v��
��
!˕���1�J�u��K(dҏh�LL�Fx�H�`liqB鲒��D E�&J�'�����j܈ �5��]��;��@��Ǳf�]���Tw˳�%ר[?�,�/n"%@�Ѻ�����ԡK���KG�����6�i!070�jV��e�������'�`-K\���uo=(H�lA����aDַ1���@ %C����n��S۷��,�w�Ɣ�%Q��؊`,!t�� (�����n�0���M$S�������bR�iaS2"�H��Z�~��{�['*r�o��*Tea5��~�:G1+�p�[����2�dO�Үv[���ۅ��9�a�.����ۥ�s}6��U ��C*�	$�RF,	�|"٘k����6�����kW�P������T˩ܘ��ꭆ�l}�w�8ʰ<q�(S.J�{��.���hA���h����65h�Zy��iDh*C6c�+��%��F����_=�RRYa<�F�+��B�@ҋ����X�X;�s<D�r��I�A�Tl�xs�V�����[�fO`݉i��;�a��|l��Z̬���sO���5gxɤd7@�x�R�F_�	V�-�Z��e�[�P�I���R�mL�+W�p�Î�(#�ŋ�h8q-��hK[�0��2g�����1۰<NuT���+l�ZO�ML��Ex=L���ݴ������8`��쁧�'גb	����Wj��l}&u�=�swk���6�=�?jT�!y�.�Şni��P�Ta��3�"94q��7ʉ�S.�L!M��57��=|�j<��U�s0�/���a��Xbރ{�tH�wJS�J,���~��ф��R$��w4n�-���!�ʝ"k�3 Od:�k�P#8�"j�J�M8�\�2�M��)4�Db��)�Y&B`&Ϯf{8��;i����8�Wo=W��·쁭ȹX�==���Lјc�&�>�;��0c8��A��l`���0`���@�w��^Ijr�.�$"���H�j>1���@��[b����E�p�ţ�-j�@��oG�/ƑJD{���S�E��#3i����_�7�eC��ă>fEʈ����PK/�	�#,7�EkA�	��1N!lf��\U�2�ʾ$Q��9�~17��B<��9��X 0���ŋ��a�L���jXy�a[|R��+I��J��Ak����7�6O.�w��$��E������Da]�r'���;��[��O�(���S�p�<\Zmbߓ}�w`�]���]���i��Jō�D߫x:K�^����V]�e	1Ϡ��d�.�{2h�5�Or"J1��U��L	Be���;��Io� /���#� "7��zg���-�#0�#3j���e�*u��i���βT'Xұ )��'ï�����~�ݺ����uO���aa��Jq#V�4�MUq��Y�*m����cj/6	��/���NȰ����ve��&���z�rDٲ|Pm&��U�쌖��d��]���H����_ۮ���� ϥk���Y���!K6�h��S_��7]���^�2s3��R�)�!�>�VN9��� u��iU)f�ȑD�\��c�=�N�ڳ4�ч1��-����S���o��y�F��/��-V�Q��W ���p� ��'�RW]'�W�M����p�K_C� �D�_��Sd}���腻Y�|L(ޛO�j��DƷ�%X��.6��|%�v�j�>/x��X=)D� a>[���a7l5�荾1l>7�l��M�3A�!h� ����-�{����� �3���|0'A����X\����[}:��flM���,Ǹor��9��'���8p�Y�7�7м��T{QO%��Zc�=����qZ��|���TH�;�!�+�_ue�4�|:0�bp���i�����u
��ghE�|)n�
.�g���hO�{���^��"�G� ���u��5���E?yoblK)YȒ�[�p��?�i-"+�ĘT~�����9�H�N��>$�:�m���\d	�|�c#_���O0ziG�yIH�u�Ύ��Fa,���֚;Z��D�+.��4�d�膑B�2�l�`~�5G�q�zw�8o��P���d�{F#�R�+c�`"�}�&=��u�E���(�:hPW��9��W�"�8��ТЄ�85�D��u_P�+9�N84^H����P�u����ē�~���_��E�I��y�����4h���8�����LxCGēU-��JQ������)��@��Q��Ӗp��Ρ4c������GW�Z�Ɣ5��l�;*[��M��]�Ys(`%?��-@#[� ��<�IJA&}:̐�/���{HT�O���9����c��hʼ]�M���	ўi�aA��3�����N �����|���^�s����GQ�+�� ǿқ2�+2����1�uc)y��Y%P�@�˱�.ba�e�fU#�X��2-�Z[�K��d���T�AF�t/G%�I-;��/Դ�����]�$���ք��2%�KC�����086��H�&SYɶ^{��~w��&�tD���>��޽���F���c�t�D�<���/<�PU�+L�TYiqg�|�����8��$ ep[��wYX��pQ^)]���7�ś�4\���Lg���mǚ�hͱM��_"��q��]����<@:g��'�4/���n��8������[�f���^���責�9�##~e?)�vܕ�*�Hp�(�~���c�G��I�T��1%�B�t�fj�Fo�\/��`"�� t�Hp��4 ZT)Wf��Q)?dt�4ƋE��w�*FhΉ;r��*�9�S�XD��>�Yk�1�,�K�p~���xd}j�fo��\�{���Z�#����S�-�|?�ue"��,z(���3CΙ��t��ߩٙ���O�]|k�i~�R�v���u�������Z	e*n꿾�R4���-���5_������x_V��O����.�.����-J�-P�Ŧ�������w����ߖ�=C�k�<%��tP�f�ϓ�ں4X��@7ۋ�|ݩJ*�	��3���6ҩ#j+��d?�kv�H�ȃ�Pyx�A��s1��i���[./�5��񞤑�S�v����٤�,!M��k�#�J��*�рFQ���hLh2	�����o����5�M�ދa��ڙ\�Bye���1���\,��� 4�f�5�9Y�Ձ6���PA��� \-��'���+��-�^�F��a� vne����Zf�c�~����d�[*w�;�v�����. _�xo!x���ƪ��:�A؉��"�߾(ƤF�I(��\Dt��DKG7�$�J��ڛF��9e��=o(d��k��\M�ŭ�\m�B� b�����-d�/�[1�.�������x��}tC��ɖ'��)�����}(�%�P����+����� ey@�nf�N���$O,~-{U*t<��[ҳ�M�d�b
p��Z���S��k$|1v!B+>&�_`eݦ�U�:c�����xg��j�L����P�PH<��IR�z�g�̐�:�	ሴ�� ��U���K1DԜC~�`�un���4�^�����;i��e��.���Վ ��=��u�
}�R��QVpۥ۰b��j���I ���V�z��Cl� �p晟A�����v�؍�[������q)v��D�K����� e�IB�ǃo������j��6�
�$�-�Ri����D¥xR�4&�I���r��g�ɗb���1U4����igs�o�Mٛ��}�@R���P�ggi�������)F���*� ��7�U�W���0R�r�����v'�����D� ������|b^&JϬ��zB���J�̊��55�ϩ`��ю�����Mɰ�cj�f�1�-�d� t�A=s���a������W�~Ma����Lh,?�7d��E j<0h���z��ŹZ2�nXżqZ��W0�J���6�	����L�t���1���gAO�G}s�8��{�J�!��=̩���J�ߏK�U��x�����l�c��֡+Gj�D��S��k!��
Bߑ���e�����Wa�~��(�o�Ȳ�؄gM�7���J~>U{���Z�.�UL�'�s/�M���0���C�='�#��:NQ�0[�4}��f5�=g�;7�ɿ�䉁VQ(��8�H݈�]�a�}�i!��(u�K4Y�{A\��ROxGuVѿE�u��6p��E�0�7�?�jN�2o�:��g�9E=h�*�>[r����6E�:���(�ִ3٘�HXKo��O�Can��0n�7ˤmP�AZD�? 5�NqO ر���R>���yY�?�Е�o���o"?hQĂ�ƌҷt�ӿ����_i���s�������%���J6-������A
j78���(�z��������u���p�)
B��e5�t��d�p�Lf�b��I�w a�3�(�Ȳ�aZ��c���og���O=X�q�ԫ;���Ac�Pk&��X;]����&/���݁��%p�k�Z�"�����eM���%�Ј[�=���*_d:�N�DZ�弦��b;wb�0��,��'k4鱘��<�F*G�r?�V��a�Z�Ls>�q݆�x�-x�+WC��F���"���Oy�ъD�]��0W����y5a 7�+29Ȏk@���g�-���x)�t��W��=�F���SoϷ]� ��pk���O��)��Fc���jzU0"3����a�va�:�c>c����4-� u�|m'�����/Ϳ8��M	YgS3�Z6����%SB�6)E��#�\mTEDy=!73#_��J�%�}9�5]��{
&0"7ڴ�&�	,����ͯ��U�Ά;q�3�س�����qb��1⎘�?�=�����sG�^��!�蓦�`��xh0�iQ�-I)���Ω�,��U����Zַ!a��5��be"'����B�Qg�"Ήo�K.@��˨�^�H|I�Ǧ��$:׏��c��s�ڢ�6>0A�A�Kr04�8�\N(����`υ��4m�&@�����M�]/QS�7���UW���$���s��˝�Ap���XQ	b'�+�/�7=v������T99x��Ż��u<#N�ou�΢�c�oQZ�ۜgg�K[J`s��H99T������+�`-_�]}��nB��e)"�D�L��cO �k0`7c�U�N�~W(��B�b)���I����¹��*e�+1 ��㟮�c0v��p;�Jҙ)�ˁE�/Q���>�8��ô(v/��]�"�߶s�2A�6�K) ܳ҉D�@�Y���:E��d�7��N�(��(��n���%�sg|N�:7�/�w�vfG:�01���R����@�����ԥBS�"G~A~�U-�HO�HeO�Y!��.�)�.�6��6��<���LG��T���/�9|��Ec3�ː��ȥ� s}/���28Ϛ���#О*i;�����Q��� MG�����J�<��/R�(!����}G�>�p䃷��LAxUI�&��q`�����=gU1������6��P�5U�U���m�i(����z����kY|F�Be� o# ~b׿]R�x_Mj&D��Ԧ��[زv�U2 �6h;T����t�W��c%�	�z�)в�ۺ�����1Mq�P��ma�Q�BDd9ޱ�gfy�-f��Q|<�fe�.<h+	���q&��
G�Ы�ZOġ��@�hW��.�E�� ����G@���%�Q*$��f��#$m[S�a����`>l@�X߷��=���I���m*mњ4I H8�
��1z�sN����ݖ�m��WN���=r�^�=	^%���W���'B�X]�;�r)`_�����wmiWs��r}ql�
�-��R#��-9"-��3�LO]�gH]]6��Q�;Q�X&6�g��GR)Dn�ZA(�y���o�Z�4-�cJ�Aj3\jg���L%3!��������c�������|�u�3���w�:�n�5���F��:tnf�o1z����+UJrbQ�B��˼���St[N�P����!�JK�,�L)X����� 
� [c}\��R��!_V��x���K��a���Rhp�s46�ʏ":����/���y�4K�l�v�3�,������"c�KR����S�)�*�̧�oɯ~$�
�1�9��%!zjI"��8Kh� �,����g�9�l���@7�$X3�|)��zM��e�ѩ�� 1��(P���܌���9�c��Y9�LZ�"���RV�� &y��`Й��S543�J�F����@}�b�,FP������4�e�z��r��J�-��²
�:������Rrb7�rM��³^%��%f��C�}:�,�9���d���]Cݣ��5��H&�`Y���Ю���!K��6����V�Y#B�-n�
������T����Yp�I*z�"�6�1���ж3x����T��~�.�oYrd<��Z��*@�7�C�sʏ:v%�U�UJ�-��1YKO�XU�D��ܹ��L����&�,;!N �ؼ��]�D��㗦�DU�1Jp�qi_�Y���?������7\y+ �ԙ�0�W�b��na4`�!�T�I���mi�[�~@��=��Y׬� ��랆�W	S�;�j�і��9TZi�8�����b$�@ ºTPJ5�Tw��Tٝ2���O�+���8k�l���7�Ƌ����_��+����	�0[�A]W��M+4`^WˀE$���M��n�b8x��	u��Y�_#�������;7�ΌVt/�QEx�Y���QV�����G�n��b4B˷{k������rT���%���,���µ �Y�m9/������e�����q��L�Nn��#]ne�lw��7bA��m*UHd�-���N<�Qp�z.��XP��������ِvziQ�66�8^ÛE��I���C(:�g�L��;RM��>$F�"c�=�d�FI���r�'UQ,{�,���Co�?(ąNr�˺
�𜚁�.���=-����$t+��l`�9��&."A�C��(FRM���$k��fy1&�B�:Nn����8�_��)>����H���9'�M�.+����Dj�(�ꦸ�6�\�Q���Z�P���7AF9���N���i�t��8o���m�lc������b 琶Q�SSjU�	�l��e��}hs8����-Q������C._�����S~��;��R���[�K
�� ��f�W���]��=����!ra�w��i�~�I_5=���#&�.�E��aQȳb���/�D�/�K� *ZSLOo�aT�5��������y�q�l;Zl
eT�B��D�"�c��fe��k���*��>}E�5�]R(�V8!�Ï9�w�VqH��"nb��S�BZK%��J���A� ����i@637i��@b���G�2����p���#�[]��RǪl�A��-�īa�"8��v�oZ���"}�u`������Z��Ò�,Q��\IGj��#��;�2������.r/@��2�PjgVv����'������"Ⱑ���HAw��m+�����R	͘L� ���ϙϋ���Ǚb���s6�Vb��q��H���G>�G�@��(�(�!������x+j��F�^ЃNQ����Ǫ���ǹ��8v��R�X^��:-���R��KZ-�-��D^̂��������X�	%�
�HB���(�sz����n����/p�z	�?��B*��f��_mb��7O��a=��N0Уif��N��D�q���;r=E[k �Ev]3�Wx���5*����Xڊ��x8���F�g�_U�ٸNg��w�wC4� �h�{l�Uȑ��!��~%�e�?8����o�O?���Gw5��"�@<2e3(U���s'+���.c����
`CrV��oh��Ь8pa�Z���B*>�k�V�V�]�_�%��?_#�����O��B���:�����2��G�Z~�������&Y�Z8䲡���'a���skN���o��="���E�n�2�1�/A����2A�L	�� �V�8F&�ٱ�=-���PϷe ���	�ʄ�L��W�L�}=�v�'L�%���%�q	;d��b�1�b�?���bj�#IX�h��\���a�&�9�l���*Π�r"�\k��%���U��P��� ��o�f�B����ɛ�S�!{D�LP�x�;�_�����yA^�*}8�$r�1�1�R-e��0{Z����Cx����G_8h|]��(.�qK��X,�k�i�*�<��NP^���[�1NxY�x\�UZA��HzܪBV�^C���k�w�eXEo�gc������Ļ�K#!���G��V�E�Q:E�d����J������y�&L�����[fL8����Z���)f���(٠RUahS��k����SFĊ���R,��*I�sӧ�n�M#3���fL��=s�P���[��r��Ū9���޼{S�!(�&q@L��֐�F�y!a�n��}��q�����(64^��Q��)�8��g�mq�C�l.�p�u���V�<sfX4�Bt�[��4�o�"�Cs-��
� e�����{���Н�Ќ>������Ԑ�[�K+gc/3UadȚ�!�u
�ب�inA|�8������u$#P�d�J�N��4�0vУ�a]�ƻ�=_�B���K����&���U����o~m3b� �>S��k�9R<5������g򭏎��!���j����:�bMQ,��s2�wٸF���+�P��|�,*/��H��c�k<In��<���N��1�9��L(bJ*�ժ����g�'g	�:4����x�_P��'^O�r�8�	TyLy����kC���U���& �c�XR�%g^��/����}���Xh�	�%��^�C+9�,J���[�oW� 
o����n�x���^��`�-�2!p�ꡪ���L�v"f�	��p��܁�E�>{�5�I�����u~ؖ¹i���Y}�����5р��[tN�ǜ���I����w;]���Щ��{��h��W�m����T��e�=���_g�(�7\:[�0;�Wݟ��碟��[g�+��[��9mO?�7�jO��N�
�����I���f�9�9e���]~��3��#�4��	�cA��&�]_��~��j�I�*��õ�G=�L �~y>罧��S��	zÙD�}<�
4Dy)��.8O�G
�����{�ʙX.�ND=&��9�'VÉ<t�����`���y�F�_��ߟE%SWg/a	�5	���&�;�jv�����1�s��zu?W��7oǌ\;�v�����gɚ�R���+*��^ド��i�5�� p�P��Vr�F��#�Ƌ��Ӌ���Xbt�"! �Do'p���SkG�S����{�N0��1��g��L$M�#	�.=�"uu[�Y�	j=_��frǠ;�2�>��g�5�e��24���
�O���%R����eȄ��o���}  M���#S�5;m��n���,k�9��j�SKK���AH�d2��=�O�u�W�֝�����Ky��K3-+�+u�>�t��_H��n��U�?|:I� ���<-�|<��+AǊb��%�L��2���<}�Z�n�_���@LS�R�G��֬ƙ�w�����d�o\��`�"ל����ؖ{S�U�"�b��S�q��ݍ�v���. �p͜x|��r��/Ȟ�@2��'o����b����X�Q��R������m7�0�~)�ﳽw��~�G5�F�L�44�-�<�ezl��AV"�v0"h�����/���u��Ԓӓg�6�� ��	T*A�	O���\�%~�\,��8���;����t�� �[��P���@�����&I^/�c�X�ex.��p������^��g��݁�b�H�'�2*v�'��]Ү39U�GwE���>�B����\���T�{�k���~@� j��C����s�MF�4h�\�{��1!�\0�^�3@�
E�{�+0�b�z��c�hX��0��H@_e#(I f���ԢM+0�4R4:S:����"|����%���f��������{d�k�,R��f�%w�T6.�aHfCE���5��)�Ba!�ym'�^�$j����y�6_��K2!��9�Dxp��`�A����oۄ��D@�nbj���ϻ�d#oK ��]  �ޣ.���Jv!ߩ���<]�\��E��1.��ɵ3����^̚Ϩ>uE A�:�y����ML�㇍���q%(ɐ�d��&���U4�A��T�m�q�	��g}"DÚ�C]��aO��&�K����������&�Ԑ�`
��@o�������}���|�_�Ȼ��?K@�{T�)�!��ݰz`M\��g�_(�w��0?�M�@�^��ɦ��.~/�'#,�B�	�>���yz�2JvOy�6��	�����Sʫ�¼�e������o������th���uC��аj�Y
�_��5���?�%�6�6�6�9\��A^�a���N�/� $i����D�{�j�Ï�]c#v$4c�ްV��O<��v�wڣT\�5�����㿘n�7�f�1� |��;�����b�B�I��$����5�/��
��	�%zn7�;��yH���C6 X�p�3Þ�
���:��"R,;��xL��������0��B�,�Ym��� F��!�@^�{��ݘ�Qe��+��Qv��}!� r\}�Q���k}y�_CMp2`�U�����C�+�K�bI�xG#��$��]c��i~��)�[��T$a�u���P�:���Q��"����>�M.�!(P���}�U����uH�c��x?��j�NfF�d�*\��nGbX@%�Y1î��I�g.�ZH�+.������3���%u�t�rL��?=�0n�T+ɉ '�ݚ� ��3�"����Fj�H�,
7d��s�ٖS�q3����ޞ{���ߌn���]C1jMw��d�y�bJ�Kv"���q��0���9�w���Ϟ�On�Z��=?�е��ᵦ�)FW#�x��SA���!`���߇}�H��I�]#.� ]��o��-�w���=�w���9"0�ļ��k�(�\5��ޕ�]�)T�>
ũ�j�L�CwK�����`��;~����w�)o���&��x�muȾ�**��i����E��&,��\b
{���b�us��-���r����8��.��ӳr����	t� jZ{6?���]�
0؅y7�ʁ;�����V_@��[�L���ț��Rh��2��ѽG/��6#�GC��U�ם�t���ɒ�a~È=��I��c��6>�ߞG�Mh;�y.*�̧����E�E^fu;�5FJr�{_U3����7ح"HU ��t<�dc��z(k�j�rcق�,������q��C>n\}�L��R�ho�!l���%��ֿH|�lھ���<Z��;��q���X]�Z�:��5����N��=cD��B̚��6o�K8� 6�a9OO[��yCNDCR(=�3�ˀ�K���:�E��J�' F��~�8�(uA�3�eIK.a.>�]&�:|�����L����!xP��fp���"��dZ���T&|��{9�Cݫ���`5�5.���g����!$���rdр��yQ�����z�W�A�>бY����p���*��l� g�pFq�l�va q�צ�l}��.O'ٍ�	ui�ϸ���XU"Jn{`8t[��T6�Z��,�,pZk^������f��L�^�*-6��U	㌽зb��|l�zL.����A�Nv�1A6 ��Ƿ� 	���<�OMyY=�n�k^�wo~-�$o���Ͽ��<=���JXe��>i9w�,H��q�5�H}�a�6%0�z�Īf��۠�,ނ��j���p)ûl��*��{AȻ7(،N	B3�5���{Ѭ���9�|Y��	&P�y|�jC�Z��:���g�ŭڽa-�}�v�w=^��xc��%΅�́�Y�����&�Go"�>��>�mcQ!:���x�� ��T�8*=Z?�' �f�a#�E^4����P��S �c�[�b�PS�~{�B��P���.���MIM�ʴn�WԠ��v���Ӯ1#�U�M!��0+g��������^.1��Ӕ*�k�*'5�����N�/P�Hsy���Z�����I��s~ � ���B���Eq�����Q눰��A���8b�_�\{۔�'t��R-뗒�d�R����<Ϭ6N��_��0�K���.~�nc�<[��i��ge����n����9��;�i�,Ol�����p��O�6�K,�6mx,��PQ��H1��$ݞe=a�`� '8�g���q\��}"c�k���+��|.�XT;p��'�� E
�uv�`�=^�K�Z?Бrˈ�;7`��^����s�!���?��İ�V�ܮXzU�7�*��ARo�����s�P���7�f��E�O��u[8H���:`�=��f�!��%���!����nצ<�S�wC��]����9�ā�A�|$�Y뙁�!BK�ky�$9��w��s��z�������h�;����	�R�Aj��N� �-��ȁ�k�~+MQ2-*�-�Y �	�N���o��ڣ"<��#��睼�G�S�,�����9�Pc%�mFW�?Ⱌc����$����}+(5��yF�|��%:�}[M�,��a����b�G�I�?��	D��L"��(ۂ���u��i�p��j�@Q��������L$�����p�M� W��/��_�p5�X���\���{�+V��}ߋ����F��=��s�F<	�^�	���lko�Zv�)k����v�
�ϰ��7�ajF,�|%/��D[!�(�q4$X5"O"E����abE��[�����Ţ�4\�-è��:RO�f̊����3#���,���үq�����-���~��r��I�sr�m�)�1t	� � j��ES�m�-����O��˥�t�3�o`�XG<Zs
Ϛ�zy0���sp�Bk^���K��¦"��4��-���p�-���~���v+�wY���g�ZBLs�eqw�DV1g�D�	���
�䠵���;���#��͔���x��(Z�jwj{X��M4��97��Ll�EP�O�N��=,�D^5�~+O��yB�9�ފ��TN��Vg�KGq���b��p+�7/E�&1}/�[�7��6��d�^S�p�0!W�/������'�KR����A.����8�w�-SS�|���s8���b['���K[�c���͠ei ��fp�G5��R,�cEX���MƁ*{�S͓��x�� �/�;��8~$p#>�4S�
�%y�p�Mp��[7b�IV�d�T���vo%IY���E�ߐ������F��¥t�sّ��]tSյ��`�f�o3cs �8Ɛb9��LH;���������:g��I�F7��d�q��^%�*(��7��i]#��/j7���-~插�����g) q�!C2h��VZa�|�?�/���.��w;U�J��F��Z��+��;+(��:�;H��5ngے��R��1���R1	H�Ax�'^������ ����+�����Nt���s��N'��7�id�iC�鲓{�;�X���C�W��Xԍ~w�)�U]�x�jq�eQ�]��YYǆ<PmN����&�3jE��=E�Z*Ś�iF�V�Xߛ�g�+V�࢛$I��4(��R+��c��V�To�}Z�j9h����[�G��T���e�}몍=Iu��s��tʭ��MbuW�@8��@b8N�MD���r���+����H�`��,̝ B5�P�T�2��-��f�3$�Kc� <�m!�ʄ1"�b��٤Z4]E}��u/��lx���?]�zQV��]{F�[Ȗ��e`�l.ڭp���O>��vd'�V�p�e�}���3�&H��ʬ��']6�;�)���)lf��1���@k��+�H
�J��gw�^uc�.˖�g�a���݋}@޲'�t>/ת u{�+3�ط{o�x0W���͑̔�]���,���Ȕ�^8��G��n�s�e=�р[��?�j���S5�K�\,.�Sϗ�V��{xy���Z�A ��^��Ϯ���h�Z�����!����c������m�<*( �jH�<j�v�i`�~�.�C=oH$���Z��3�׌��>���%�}r�B?`�cQ�8�SQx<-�]u9E�<?�%'pPL!�#��.wU�B��z1tێF!qtd����B�$Խ�������{�'���Tr��6I+
����/�f֫��� �]��(��F��+@G��hh6/מ��&]��D>����/mFU%W��,f�P��!`*��9����ҙ��b��%�Pq��~}��g��b��	����>���oET%L]KPV�:s�k�j�I������V!?7����X(Z���.ͼs9?�����������p�4BLԺ�6O֪��탤�,KȜR9�$"A��$XY�Kˬ��ޛ]���ա!$�h�WC�>�(�zs�P��fFp�[�>i�9������� �2��FE��GeOO��,˓X^8N�,C��}{�h0��<!Cl=/IO�h����Sձ��琄�yrp3j=�`����=��^M��%��w�ո��,�VK���:�pc�G��1^|�8�D����<ج�K�e���l��>c�����3�NQ�C�hw��NԌ�����	�t���dld>�N.X@�.�?�H|��l;A�M�z���f�����R���'b���T�XF=ؿ&�zz��m�9��P�J|���r�0Δk�Y:��4y���*��5�7$�)�n
��b\[`P�&Ŋ�?�����p��T��n���<���Y��>[3u\���O\�|+ �H�7
Ȕ�Mv�2���j��
�5Ά JL@�@tO�m�C�;���� ���#��3_��}%���;�%�#P�P�SԔ�Lc$Ƥ��OPj��!��A�˖#=�w��R
&t���^�c�ڵ~}m�Zs�v��7c�{-�ʉ��p���#��b�I�`� �+|@LG4��}j��e$��K��K�n�89ϯ1����oFJ�a-I�c�m`�%�*-�L ��,#�:&�Ԅ(Yj����]��4���Rп��iw���JT�;��p"��[{�6
��M�z�0���:7�,`�8���\�o	^��	��D$�""�s�~�&�q�h[�/E-����)�XL��K��I��mUf��h��_݃o�$�����ٟ���u��<��!Luj�7�(h!rz��Rc{���6+�SV��0�7w�A���!L����T�?�BEL����jj=@'!߬LȔ!�5�똡���bι����R!}���lۊz����l�L�*�eh����ё��[�� �B('c�gx�xHB�ʚ�g�Nc�a,H��`�C�,�i���s���)��ek��%� �I"��c��|2�Lr
<D��o8;9{c���Ϸ ��تn\/���~e딹�u��(��t_yJ���!��*�h�>)&�<�@yX���"V���ް���޷�B)�a�`Z� K�<���.E����;" �6���;\`uՠ���u��<�cj~���1mtt��[Z��k������J'� S��ح���Y�	�ϖ �"e��9�:@˫W�_�`�� �rO��^{��G�F^IL�%��ڞ��L�+G��d�T��2}F�F5!�?T+��0zi��\�޽�3�e�HL|�FȌI��?�2��S��[�_�\>�P��5�ۘ� �E��i���e��&/���b�����AҨ�Oə�Ew���_�����{H��+ӕ��M�,�vF��t������_`t� 3ȀS��/o%\���y|J��L��!}���c_bC�s��|���p��l�{<<�v��I��@�2��;�wH
��Sb����X�2��#Bj���*������	���`��{�����1~RI>�"Q�R9n���\���}ַ�� Ô'�ՠ�n']�DQ�z���\�&CQr.?O
�?�R�aŨь��0���K�E�(%��0��q\g���P�f�h� �U��7˥�5���/�ȯ-[��RY� [.tgM��yYI�.:���Ls�g�.K��v9&�:7�X`Y�p�|eʇ�3I�D�Af��OID���Y�1���0��Q�0p�"8
��`��8�lNCT9�V�,� ��!�!ӦohHH;���_XRTw�{������E��w���^��e�մ���(H� "=G�Wn��s�|�M�"��p+܃���c���Q��b�<�(#���S���F�I�_.э��`݃ xt�XBy�g���}R-�����_����R��I��G� b 
?��Fr�ْ�b�N�9-T(��e+��|Hq�)��n����0"�o~�jUN�-���9���Z�c��^#�Y�Ư��jZ`soh;����;�:!�D�-(�XU,�\]�Iv�ZQ��hOg8�8y��~H�2"9CC��7Q��n�عk~HQ�_�z�b`�����$��e�u�P��A�[�A�����&��P2!Y�������hz�рn�J�_����X��>Rh�ImGUI��a�{���_�e�;F�N�p}�3b9��(K�5V��#%�7/"�m��B�_e�6�Xd�3���I�t�t!����c�C����4�5�X�+�V�S�$չ�� $����f����4��c@fU�l>$��?�}�������l���"E$����&��ĳZ�|_��Ņ�3A���E*Пs`k�O�N�gYJa�/.�ńa�q��f�Հ�&�}g���7�1ЪeH��n,�W�E���KP���N�@���0�8��1u�m0ڿQB��< ����#���@-e�xgS�|�R��t�;{+��m�P�㑃5$��L,.��f���rWy�n��@��
��0��O>��/�n#�F����\�� ��wTH�qD0�u�	��4s���ʚ� QYB�m-�Aޑ���_�Y@�C�y9���kw��6���4K���c|����;�)�TM鳦�S'i*��g�d�q7sazB���t�x䏗�(9%_�_��fNA¾GD��ѐU4A2w`T���#� ����po�3�ͨN�����!'u�,{�Z��wf����.y�؎l��M1��Z1p�&,�N�B���ߖ���P�ȗ�T3,����c2lZ��K���Z1�{�ǖ�y.��ҭR�֊�\��I�-���!�{�A���2�}P�1�"�O+A?
�S]_K�o���R�}���m�5&o^L~v�#�{C}�bB�6j��iB����(�(_x�E{[ʚ��eN�P͈�ǧ��77����+��f�hS��������[S�9��<� Q5����侯`i��k�S��� F�<)����V�S(��QUٗ�>���M�(�I���C����:k$�v6�ƅB��������8Z�������u("<��x��~��Z$�s�Nz ܃���"|���Ƭ�?=�`�A0t����;���.(0�w�֟������v�;
��+)Oy�������t��{��pQ�����J�FSФ���"���XX���R8D�c�	o���|G;�'<*�Ț�F�+�2�z�ƋVC�}ir|�C�N�98Z�M-%�u�P-3�qz�敖�����͍<�1tھ��0)�����Ɇ@㫷OJP��iux��_�q㚆����О��}2Ȳ|��o�2���K�$8&O4��=���)��a�yP-%]��g=�3��� �ĭ��!{�#	����Ԣ�gĄ3 V��O�;�|�l�� �>�9Џ��ai���J�p��J�V6�E4�.��������~���|<��r}�<;-{/gj���a\���` Bn�����?oD�-S~&ܺ%4�z���Hݹu1�z�g0�=o��>�q���)d�#�9��(�J�ˬ��BU�2r�Q�e}���"Z�<^^D���)���J0IV��1�Թ+�bK3o�1̾��$h��\1���m0�q���r�f�l�۠��Դ:28MPx�@��J2ePa�U�P��HȺ�(."��h&Ɇ�K@e´ʾ�旾�u\��Z��� �r��A��/���S����Q��{���\�`��[�74��6��|כ�$=��`���&�w�:�9p�}����́�1[P��T�d/40�+db��j*Qp[Al��6ނ������s��~��|f�?�소�7S��1��îNv�}�CPA8�7���BF��7I-�~f&֣��<@h�}?,�TD�c�n�r^c��)(1y{:��Dl���>Jȇ�p�Z�p�'vmI��4.���G�:�iυ4�O�)�K����Iq�1��^���Og�W�(���&`UFaX�����Dj�r_A��Ce��U &�,��>��L2���:L�'PX�#�l�a�D��"�����.��<��	��2�?��.�߶��(޶N|�FD�t�Om�J9��ۜ�D`d�K�jz�鴔�������b'M�Q�#%u}N��'��!A�6�[���<F�+������p٭E������Vu�NQ�~*8�(e&��B���,|�r��J�`@5b�YS�:�0�(����̓�;�;��nǾR<Y�N�'f@a��C� P��}i��c���z)H>l���,��H
��%[Kj�5չ�ԤbFB�k���7!������(h�o�y4����-��Y��X,������*��^����~GkO�%<�8M���R��������Bj�\N��N.�;N�[R��rCԊ�A�2{���c89>�K��K��B�[��p�g���tu��(�}�����8���rzw�Ѫ?�=,&qx=�H� j��٢�	�:��-���憼z0�t�Qa}���_#CpJ����B����F�� �*�����?��$�el�	J]��Ud,�r5�������1����;wE��W8��ru�;>yoL�>I�q\L�����;�jڋ׽(�:5tNOW���0lL]H���٨u�ì�nYr����"�S+�h��H�����Ȥ�*��m�F���F
�fC��Ɨz-0�<t������P�k Q�r[���Cj���X�ޱ�������њp�� 	i�y�@��5J�Ո�'������3�F@�4�D��bX_�vS��R�p[����J���V�[ ?S���Y<7?�� ���R������3�ph���SsP��Hu�/��\.��,*�\s���Da��B״H�E�T���(�qAx�N�!s<0Y�Be�2�O'�@ i6%�G{�Z;d�.�Aͯ'���#��I�B�}��F�b
 ���7p
��Y���4�t��.
/t�OVmbG���K�ߒ�.ZJ��$��{�f\�TbJ�$)�<Qw^�M���������=&�`�=ث0,�*D��c�
f���*����*�!���u�G�JG�溗\"�ǳ����U�O\��
���M��m	�H'4�f�����R"�v��kr���
rB5#q�v3D����}���]�?�|��j��6J��H�r��_oGO"��U���j���W3�Cu�:����<??�~����~�/��R ��7= 04N���k6ݽ���;��#�Y����z�2�qQb#�
�ɱ������Vv*� y��0\��]����2��_�bo�r9d�b�6��������s��,?�lZ�_�	x�)1IǠ���٨�#wi��cn�6�m�0�'�ܞ��sj`�V{C�T�þF��ۦX�H�tf���!�Ysk�c��^���J9�� uI�0B�P�%���p0;�U�d�~�ˉ�f���?'�)Q����&.��ѹ�G�_.�8}��DV����ը&F,�2C���dzdrjE��������}��Ӎ�9z�|����#Ȥy�v+�Fg@S�� �`������~ngߊsve=�턑�W�ZQ}<#��"kv	����H�K��m����@�2ͨ����{W�\똡�~�we�ljx�/z��uK�C�����H��ڪ������B���/�;�U�,T��']m�**/�(u4���1i��k�Dr�덙{�C�Bx:j���` ޵�b;�ebZ˽%�<#�MnPF>*roߎ1W�F�Y�ɗ�eԶ�!R�\���1S<����~��i��o�Š�@IO�(��3�G-ň�t�j���f#��ך���������SfP�o�BZ=�v40^&r?�ͩ���1KiZA�,����p��T��a���I J׶$��)������ICϹ��F"�C�`��K5|$��l�驚�o����o��4�H�Qa�P����Oq��v��FfpH�,@���>�wWa��;$�n�h�O�}y"%�L-���ͿOs9 �� wm35"�ݏ�L������2��=E�h[�^B��3xUWY�-�I,X�6X��*�
%�6!�^.x��4ۮ��N����5;T}���qj����Q�C�d���x�E�Ӄ�L1�W?g��� kU=>�o%�(n�/L7�� ��I�R�=�t�1�v�A��C�mQ'i�ɞ���f��6�#�p��p�b��;`�:��ˣ�(��\�����:�T�T���M�q�P�v&Z������9�D�i�(�i�M����5mJ��1����T����"`�6F����q�C�_��{�^�U5�5��+�����Q����CZ"�:53��|����u���D���W��J��+�;���X��nQ$��ӑ4�k��Ɇ��`�x"��j��ҽ��H{a�<���j��"��{�'��q�l�Q)�26��=��_m�A Ԯ����	3i�8t�˱ Ð  {����čA�[���aM�@$�q˰I����ޖ���K1u��~�+c��L�X"���zWX�Z��j�b�ݤ�"�4�Х �)��F{�k�Y(u/x\�5������~\���F�i>�������!]ךwE-�+ga~ǫ��Aڗuz���u���-D��I������t,��i~��2Κ�����55�h�՜2�?;<
���e~O�[��V^#�vP��ۥ��A9.���5&���`h笴Jj��$(�����ПJ;^��I��" �QI���>���VF�Қ�-������!�J�*������\"l�e�u����Q�|sN�����K7f��{��Qܝv�(��S�z��	-L�:1f� �����͔�q<=��OfK��w3#yƦд�%��W��:j�F2��ʳ��~�
P
�<5�]ׅ}��
���j7��d�U�]�rj�*�E{B6�����aѫOF��M��rB3���w�7V�U�Z�������u���9㠎?8�!���	n�U�~z����Fzzk�^z���~����9s�}%0_l�1����U�dG���q��F����X(�	��=�%Բ!b$�E�@�`��E4���ܾ���&�s��%c®c��H�w"hD>,{���ۣs��m��^��pG7ނ�D:Q��n������./�7M�'��8R���w�!7�N-��Q���3��t\���\�n⡈���ߤH%�4�N����$-7�oK�$t�whd �M	g!i44M���Ꞡ� q�w
��
�K�,͵r��]�v��z��,�`	ʁ[�q��9�N�F��H/�� �'V�a���:2)5΁��k Q��R�	t�E��B� ��gc���������u.luDu�Y����
�]+bME[Ȓ��I�**�wc��<3��cz�n-���� ���/5�U=Z�����b���(�1rOHD�rG\(܆��-+��<ּh��u�2�o��b<79��ۈ{�@����]�Kp�C#-�41�n G��>Pa)+L������g�h@8��0���ǜ����M�"i7�j��;y: )m��ӧO9	%�ٹ�靣�����>�����(���a��A����x{�q�i�֗:`�_���8 ��:oܙ�܎[����C֣�����V2�6WmK�8���?Q|�>4�$�M�b�1>%���.K��ƖR���8�9���Fz��5\��NP��X�FR32ňS���}WU�tE��D�C� �_��;�N�C�lU�M;�e:��ܶ&,XDY�zܠ��p�'��nx�r�����Y	�ۉDf���]���A����|%�H�f�N��t�Y0&��Z����c&���?0�6yf:ͭL%3e*Ek˽�(PEL}��6.��Ō��++�,�d : '��<�Ԣ�:��i�t����K�X}�����;c�4x�n�����r��L|�0��M�>\�޶{��e��3�C_]jP�����H���9�D%�t�9Yaݙ��}�g�?�����ty3������u�h!�w;Am#Nd�u��Q�ڋ/�qG�V0ޮ6w-�+��j�/A@#���IhuBJ)�q�5-��*S;��=J��؍���}�����L�7����db����y��M �!Ih� �>����v�N�:� ��<w,�F�l �Vd�:�Y�6lɚ��z��@Vw��l�ƚ۱w��}�܉O����2�hT[�)�*2��R���c>��r����F6�4�T�^���^�Ag%���8Yj�mؠw���9P��U�r��zeM������>$�_��?{-�#m�xX�ӭ���Ҽ�5\���b���1����_������/�%y{���pFyQ�ѡ;m}�-H�F1���Mz�^Y�m�~L���=�@U7'��[e"�Yj��A�$FZ�%V��VP�h�4I/`̂,6�ɚf�N�����`D@�"!B�,r�/&�l�VY ���I*J�}�^��.C�!.�n�=��~�\�<��:�2�p�M�{��A��1�����S��](
�6\�����U%8�>^ۘd�7*�#&�N�9�DT�fKq���%�	�8�}����M��(؛����r���>����9�_�ܛ-KEW���k��k&�f���-�L�(���\@3���>����:�ΞY�H��]_H�(i�$�u���H����+<��dN�l���K��%[]fս"B��1�v�`RUS^�%-�X̥�yg�)=	֨�
\_(:�(�>�۶��)o�l������b]Tļ�d�X��Kwb'�v��|.�P���ŏ���gZZh�k,�Ʋ��n�LSzy"|�n���?��]s���02�Zr��u*\�@X,k��vz	������̩/ �✘�M�k�st�j��V)!���	y|Lwv�,�t��V�	&-z�ؙ0��5#���C`+ 7�.b�@�4C/���n�"d�J�Ik��!�/Fe�C�˪"❂���iT(o�.�'r�uB�����xg�
_� �(�]3�V�8h��Q{�F�ԫ&d���Pu��@��
B+�&l�ł� ^z��(딿�<]��m��XŔ�!��/l��)��#��"� ���s�POЮ��1ǎ<�� ����&��lf���o�eY]ɦӧ�o�z�@��S�e�[�q N�S9,����*8D��V�_��ۿ�zR� TF���R��0�.�ymi4=`�F�ǗG���+�����E���H�t(8����EbHt���X��>���怨/?�[��cIr��2����-s	��V�y�nM#}�kM�Ә�(�C����.��z��6�`]�龏 ��:�`��FDD��������JN��*�M�#!���5GvaH��)���7��v�m1�����'��,}ꪜ|Yd�����~JP���K� �$�6H��Ǚ��((�mH�&�2��E�8<�Z����:�e�]��
�j��"�5�0M��i�3P��T��C�I,M�_�L��7�� ��~+��A�n_��K�L~N�-X�*�V8������QR�)K�C��V~eD~6(0+�EH�g���g.��<_L�lF-`#3\�	���`�/�huE\��!���^�w��ള�6�g�4_����K&��2��og�z]�h���#����ѱT���L���,�[K�I�� R�m��W�p#�Yq�!�"��:Sa�c#kZYP`̹RzZ§��;�C���i��9jK�lp-�9��K����<�t������2�}ê�O쌀���$X�{���� t>r�0� �ށ dN�w���HFsI�'9l~E��2kMK�"�kI�ܱ�r�6MW�w�ˋD1@��d�����b��};}r�.2���a�~sD6��[$e���qx�yޜ72����Z��f���(��Q&0)�����c��|~Vu�t[�:�'�rH� ���gю1���fK���o�3V�n3�	���0��c�I q­]J���|ۦ�ږd���:Ñ�i�����ݨ��ّ��hP����8��4���]�qU�sF��w��W�[Ā��#���,����4r�:�Yw@c?�q�K7P^x��OE� ̵%�R��9��i��\d�-��cOC����!�V���������=v
�Q>�v��|Q�����m�W�P��l	�Dq"<�EI�-M^��.-)@�z���^4]����'}%��S|T�-��1\�Q~&!-�H��_��-Q�Ѡ �����%o�����M/%�����ɤ�21r�_�F{�*��6v�p58���ZG���7��֒���[�)-���zN�L���},c���ye�l�s�^�A����/����T���ID#��"ZͿ����|2�wȖ �ՊR�p��fف���7�������+;r�_��*$;b-A����U����$�D�T�w�9��;�b����[q��j斉�s��@l�Ax��zx�6���Q#H�A�ҸO~�5��d���cطp�¤�y{K�8˄r�!�P%7�9kKr���j`d�Il�5_>�%��Z�3e�H�_�|\?&�"�,A�o�$��d�a��u�9��+k�P-���?$� ���ר�}ӱB��@Ō"��+V1@����e ��A����:�+�����^�O��!uk��ȭX�YLy�!;]�R��{����^f}[W�,���՘n1s�����y��Q�f4R�f�4��s��@���ޜS�A��af�Sޤ�H�.�)t˖�67���@��v��VBA�Gs{U�&C����ct��\?��A6F����҈W��gSGy+d%|�d��(3�vm�1�������^F�l�w³�'*B�����,���i~_>�R	���}9��ik!H�t韬/A�u��tC��D����N­����m���Inz��� ��/���� ^}F�u�],`L�lU)4��
�j����m`�����@������q�������	҃~G�E�6͸�	�?#��	r��W�1��Qlt�|��x������{ׂ��}�k"i�g�������O\i*�';ڒU�A���M��#GJ����C��xk��8�f�N�Jp����N[&������@f���a���DP#�A�󘰐��u�V� �P�f�-$�*;ޒƊw������Oatϕ�vz���g��<{��8X�Pf�tQ�ꉕ�%�6��!��lfW�H���O<�
�K�㋽:P���E���wb"N�`��V��)9!��)���	G�y�X@ym�	f��s.0GJc��eI;S�
��b��3����鳓�Dc��sw�A����Jom�k� !��G�FNNɯ4�{�u�#L���3(Ȇm��&l@/�W0�������祶J㼯#Q���`�R���4B��w��X��q�{'�H"8D˿\��9Zr�
@ͪY�֧x>Ԡ�8��ĞX�1蝸�'>�aneXS$ㄐ5�|L8M�]���_a��p}4�s�U*3�>B-� �u�����.��Wr������-/����DG� r�ۋ��si�qrS/P@��he7�$����x���3֦d�fmR/�V{#h$��|~ab�{i\���\��z��� �~�!�f��A�2��	Pe�ɗ~1��(q�0�<-ƥ�M�;9>�����X�8AXn���ṻ�ڝ�/�'O�L����E��o��3���)=�S�	
0 �i#�b���%�8{�|�v&����9䠦Wz��}h�6(�;��Y�C5�H��T��V�h­�N9�y16v5��p���u���ջf�Ix���|+�MMQ�:��M�T��1^]�0�'��O��q{ۺ��cp�}/�S��@3v�ɓ:�r��q�50�'n�����	Ŗ�S!y~�F8�����ڽ(�t����D����d��O��h�>�w�(��>AG�����^� K��<^�k4�Rʩ�o�����9�?�) �ί�Y�K)�t��]�l�'9�f��H���6 ���x0�Q�ǆ-Yo`��Ę����	~ ���G��H$Ɏ0�N��D";u�r�I���u!�Ca��+`�biz'
�f���h�-���e���N�$����צ��VIM��4�������}�X��iH6��g��@�RS8���I��"�"m�m%:�x���:a���A6�d�5���嚑��q�wM/O�f0&��0�9�4�� ����i��m�s];�BI��~��0�c'w�4?�V|��Y`z�D���}���B�fM� Ks�>��X���K=�H�'Y<�U	��>nL@�W쌓��=���Z���b�u+>��Q�/hQ:��nf����ϲ�.%�����P���u��^��Av��G֖���_���������kN�&"$�q��7U��`a�Ř�^Ba6�Y��[�[��p�!~0豀��9�">M���cyQԮ�/��N��i9i���Q�)�K�8&����SC����x�Պ��'W�$|�¬2�٦[��*	Lٮ�Tf�4B�A��U���S��24����nU�x'��L�'C��G5T�'M�=$�:��5���I>|���a�i Oa������>R�Fݰ��-�咄�"��&�z*h���<���H��LKpT�g�kMO�*(�<T-�M�\�s���.�肟V2�������Ҙ