// soc_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,        //         alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,       //                                    .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,      //                                    .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid,  //                                    .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,     //                                    .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,     //                                    .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,          //                                    .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,          //                                    .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,          //                                    .vid_v
		input  wire        clk_clk,                                    //                                 clk.clk
		output wire        clock_bridge_148_5_out_clk_clk,             //          clock_bridge_148_5_out_clk.clk
		output wire        hps_0_h2f_reset_reset_n,                    //                     hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,      //                        hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,        //                                    .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,        //                                    .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,        //                                    .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,        //                                    .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,        //                                    .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,        //                                    .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,         //                                    .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,      //                                    .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,      //                                    .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,      //                                    .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,        //                                    .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,        //                                    .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,        //                                    .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,          //                                    .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,          //                                    .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,          //                                    .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,          //                                    .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,          //                                    .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,          //                                    .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,          //                                    .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,           //                                    .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,           //                                    .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,          //                                    .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,           //                                    .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,           //                                    .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,           //                                    .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,           //                                    .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,           //                                    .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,           //                                    .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,           //                                    .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,           //                                    .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,           //                                    .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,           //                                    .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,          //                                    .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,          //                                    .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,          //                                    .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,          //                                    .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,         //                                    .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,        //                                    .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,        //                                    .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,         //                                    .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,          //                                    .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,          //                                    .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,          //                                    .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,          //                                    .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,          //                                    .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,          //                                    .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,       //                                    .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,       //                                    .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,       //                                    .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,       //                                    .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,       //                                    .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,       //                                    .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,       //                                    .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,       //                                    .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                               //                              memory.mem_a
		output wire [2:0]  memory_mem_ba,                              //                                    .mem_ba
		output wire        memory_mem_ck,                              //                                    .mem_ck
		output wire        memory_mem_ck_n,                            //                                    .mem_ck_n
		output wire        memory_mem_cke,                             //                                    .mem_cke
		output wire        memory_mem_cs_n,                            //                                    .mem_cs_n
		output wire        memory_mem_ras_n,                           //                                    .mem_ras_n
		output wire        memory_mem_cas_n,                           //                                    .mem_cas_n
		output wire        memory_mem_we_n,                            //                                    .mem_we_n
		output wire        memory_mem_reset_n,                         //                                    .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                              //                                    .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                             //                                    .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                           //                                    .mem_dqs_n
		output wire        memory_mem_odt,                             //                                    .mem_odt
		output wire [3:0]  memory_mem_dm,                              //                                    .mem_dm
		input  wire        memory_oct_rzqin,                           //                                    .oct_rzqin
		input  wire        pio_chaos_done_external_connection_export,  //  pio_chaos_done_external_connection.export
		output wire        pio_chaos_reset_external_connection_export, // pio_chaos_reset_external_connection.export
		output wire [31:0] pio_chaos_shift_external_connection_export, // pio_chaos_shift_external_connection.export
		output wire        pio_chaos_step_external_connection_export,  //  pio_chaos_step_external_connection.export
		input  wire [12:0] pio_chaos_temp_external_connection_export,  //  pio_chaos_temp_external_connection.export
		input  wire [31:0] pio_chaos_w_external_connection_export,     //     pio_chaos_w_external_connection.export
		input  wire [31:0] pio_chaos_x_external_connection_export,     //     pio_chaos_x_external_connection.export
		input  wire [31:0] pio_chaos_y_external_connection_export,     //     pio_chaos_y_external_connection.export
		input  wire [31:0] pio_chaos_z_external_connection_export,     //     pio_chaos_z_external_connection.export
		input  wire        reset_reset_n,                              //                               reset.reset_n
		output wire        sdram_clk_clk,                              //                           sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                            //                          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                              //                                    .ba
		output wire        sdram_wire_cas_n,                           //                                    .cas_n
		output wire        sdram_wire_cke,                             //                                    .cke
		output wire        sdram_wire_cs_n,                            //                                    .cs_n
		inout  wire [15:0] sdram_wire_dq,                              //                                    .dq
		output wire [1:0]  sdram_wire_dqm,                             //                                    .dqm
		output wire        sdram_wire_ras_n,                           //                                    .ras_n
		output wire        sdram_wire_we_n                             //                                    .we_n
	);

	wire          alt_vip_vfr_0_avalon_streaming_source_valid;            // alt_vip_vfr_0:dout_valid -> alt_vip_mix_0:din_2_valid
	wire   [23:0] alt_vip_vfr_0_avalon_streaming_source_data;             // alt_vip_vfr_0:dout_data -> alt_vip_mix_0:din_2_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;            // alt_vip_mix_0:din_2_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;    // alt_vip_vfr_0:dout_startofpacket -> alt_vip_mix_0:din_2_startofpacket
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;      // alt_vip_vfr_0:dout_endofpacket -> alt_vip_mix_0:din_2_endofpacket
	wire          alt_vip_mix_0_dout_valid;                               // alt_vip_mix_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [23:0] alt_vip_mix_0_dout_data;                                // alt_vip_mix_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_mix_0_dout_ready;                               // alt_vip_itc_0:is_ready -> alt_vip_mix_0:dout_ready
	wire          alt_vip_mix_0_dout_startofpacket;                       // alt_vip_mix_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_mix_0_dout_endofpacket;                         // alt_vip_mix_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          alt_vip_tpg_0_dout_valid;                               // alt_vip_tpg_0:dout_valid -> alt_vip_mix_0:din_0_valid
	wire   [23:0] alt_vip_tpg_0_dout_data;                                // alt_vip_tpg_0:dout_data -> alt_vip_mix_0:din_0_data
	wire          alt_vip_tpg_0_dout_ready;                               // alt_vip_mix_0:din_0_ready -> alt_vip_tpg_0:dout_ready
	wire          alt_vip_tpg_0_dout_startofpacket;                       // alt_vip_tpg_0:dout_startofpacket -> alt_vip_mix_0:din_0_startofpacket
	wire          alt_vip_tpg_0_dout_endofpacket;                         // alt_vip_tpg_0:dout_endofpacket -> alt_vip_mix_0:din_0_endofpacket
	wire          timing_adapter_0_out_valid;                             // timing_adapter_0:out_valid -> alt_vip_mix_0:din_1_valid
	wire   [23:0] timing_adapter_0_out_data;                              // timing_adapter_0:out_data -> alt_vip_mix_0:din_1_data
	wire          timing_adapter_0_out_ready;                             // alt_vip_mix_0:din_1_ready -> timing_adapter_0:out_ready
	wire          timing_adapter_0_out_startofpacket;                     // timing_adapter_0:out_startofpacket -> alt_vip_mix_0:din_1_startofpacket
	wire          timing_adapter_0_out_endofpacket;                       // timing_adapter_0:out_endofpacket -> alt_vip_mix_0:din_1_endofpacket
	wire          pll_sdram_outclk1_clk;                                  // pll_sdram:outclk_1 -> [alt_vip_vfr_0:master_clock, hps_0:h2f_axi_clk, mm_interconnect_0:pll_sdram_outclk1_clk, rst_controller_001:clk, rst_controller_003:clk, sdram:clk]
	wire          pll_stream_outclk1_clk;                                 // pll_stream:outclk_1 -> [LOG_Generate_0:clock, alt_vip_itc_0:is_clk, alt_vip_mix_0:clock, alt_vip_tpg_0:clock, alt_vip_vfr_0:clock, avalon_st_adapter:in_clk_0_clk, mm_interconnect_1:pll_stream_outclk1_clk, rst_controller:clk, timing_adapter_0:clk]
	wire   [31:0] alt_vip_vfr_0_avalon_master_readdata;                   // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                    // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire          alt_vip_vfr_0_avalon_master_read;                       // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;              // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire    [6:0] alt_vip_vfr_0_avalon_master_burstcount;                 // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire    [1:0] hps_0_h2f_axi_master_awburst;                           // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                             // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                             // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                            // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                               // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                            // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                             // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                               // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                           // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                            // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                            // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                            // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                            // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                             // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                           // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                           // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                              // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                            // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                            // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                            // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                             // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                           // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                             // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                           // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                           // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                            // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                            // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                             // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                             // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                             // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                              // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                               // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                            // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                            // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                           // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                            // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          mm_interconnect_0_sdram_s1_chipselect;                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire   [15:0] mm_interconnect_0_sdram_s1_readdata;                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire          mm_interconnect_0_sdram_s1_waitrequest;                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_0_sdram_s1_address;                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_0_sdram_s1_read;                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire    [1:0] mm_interconnect_0_sdram_s1_byteenable;                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_0_sdram_s1_readdatavalid;               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire          mm_interconnect_0_sdram_s1_write;                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire   [15:0] mm_interconnect_0_sdram_s1_writedata;                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                        // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                          // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                          // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                         // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                          // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                            // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                        // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                         // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                         // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                         // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                         // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                          // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                        // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                        // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                           // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                         // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                         // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                         // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                        // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                         // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                         // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                          // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                          // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                           // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                         // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                        // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata;  // alt_vip_vfr_0:slave_readdata -> mm_interconnect_1:alt_vip_vfr_0_avalon_slave_readdata
	wire    [4:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address;   // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire          mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read;      // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire          mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write;     // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata; // mm_interconnect_1:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire          mm_interconnect_1_alt_vip_mix_0_control_chipselect;     // mm_interconnect_1:alt_vip_mix_0_control_chipselect -> alt_vip_mix_0:control_av_chipselect
	wire   [15:0] mm_interconnect_1_alt_vip_mix_0_control_readdata;       // alt_vip_mix_0:control_av_readdata -> mm_interconnect_1:alt_vip_mix_0_control_readdata
	wire    [5:0] mm_interconnect_1_alt_vip_mix_0_control_address;        // mm_interconnect_1:alt_vip_mix_0_control_address -> alt_vip_mix_0:control_av_address
	wire          mm_interconnect_1_alt_vip_mix_0_control_write;          // mm_interconnect_1:alt_vip_mix_0_control_write -> alt_vip_mix_0:control_av_write
	wire   [15:0] mm_interconnect_1_alt_vip_mix_0_control_writedata;      // mm_interconnect_1:alt_vip_mix_0_control_writedata -> alt_vip_mix_0:control_av_writedata
	wire   [31:0] mm_interconnect_1_pio_chaos_done_s1_readdata;           // pio_chaos_done:readdata -> mm_interconnect_1:pio_chaos_done_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_done_s1_address;            // mm_interconnect_1:pio_chaos_done_s1_address -> pio_chaos_done:address
	wire          mm_interconnect_1_pio_chaos_reset_s1_chipselect;        // mm_interconnect_1:pio_chaos_reset_s1_chipselect -> pio_chaos_reset:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_reset_s1_readdata;          // pio_chaos_reset:readdata -> mm_interconnect_1:pio_chaos_reset_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_reset_s1_address;           // mm_interconnect_1:pio_chaos_reset_s1_address -> pio_chaos_reset:address
	wire          mm_interconnect_1_pio_chaos_reset_s1_write;             // mm_interconnect_1:pio_chaos_reset_s1_write -> pio_chaos_reset:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_reset_s1_writedata;         // mm_interconnect_1:pio_chaos_reset_s1_writedata -> pio_chaos_reset:writedata
	wire          mm_interconnect_1_pio_chaos_shift_s1_chipselect;        // mm_interconnect_1:pio_chaos_shift_s1_chipselect -> pio_chaos_shift:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_shift_s1_readdata;          // pio_chaos_shift:readdata -> mm_interconnect_1:pio_chaos_shift_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_shift_s1_address;           // mm_interconnect_1:pio_chaos_shift_s1_address -> pio_chaos_shift:address
	wire          mm_interconnect_1_pio_chaos_shift_s1_write;             // mm_interconnect_1:pio_chaos_shift_s1_write -> pio_chaos_shift:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_shift_s1_writedata;         // mm_interconnect_1:pio_chaos_shift_s1_writedata -> pio_chaos_shift:writedata
	wire          mm_interconnect_1_pio_chaos_step_s1_chipselect;         // mm_interconnect_1:pio_chaos_step_s1_chipselect -> pio_chaos_step:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_step_s1_readdata;           // pio_chaos_step:readdata -> mm_interconnect_1:pio_chaos_step_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_step_s1_address;            // mm_interconnect_1:pio_chaos_step_s1_address -> pio_chaos_step:address
	wire          mm_interconnect_1_pio_chaos_step_s1_write;              // mm_interconnect_1:pio_chaos_step_s1_write -> pio_chaos_step:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_step_s1_writedata;          // mm_interconnect_1:pio_chaos_step_s1_writedata -> pio_chaos_step:writedata
	wire          mm_interconnect_1_pio_chaos_w_s1_chipselect;            // mm_interconnect_1:pio_chaos_w_s1_chipselect -> pio_chaos_w:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_w_s1_readdata;              // pio_chaos_w:readdata -> mm_interconnect_1:pio_chaos_w_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_w_s1_address;               // mm_interconnect_1:pio_chaos_w_s1_address -> pio_chaos_w:address
	wire          mm_interconnect_1_pio_chaos_w_s1_write;                 // mm_interconnect_1:pio_chaos_w_s1_write -> pio_chaos_w:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_w_s1_writedata;             // mm_interconnect_1:pio_chaos_w_s1_writedata -> pio_chaos_w:writedata
	wire          mm_interconnect_1_pio_chaos_x_s1_chipselect;            // mm_interconnect_1:pio_chaos_x_s1_chipselect -> pio_chaos_x:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_x_s1_readdata;              // pio_chaos_x:readdata -> mm_interconnect_1:pio_chaos_x_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_x_s1_address;               // mm_interconnect_1:pio_chaos_x_s1_address -> pio_chaos_x:address
	wire          mm_interconnect_1_pio_chaos_x_s1_write;                 // mm_interconnect_1:pio_chaos_x_s1_write -> pio_chaos_x:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_x_s1_writedata;             // mm_interconnect_1:pio_chaos_x_s1_writedata -> pio_chaos_x:writedata
	wire          mm_interconnect_1_pio_chaos_y_s1_chipselect;            // mm_interconnect_1:pio_chaos_y_s1_chipselect -> pio_chaos_y:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_y_s1_readdata;              // pio_chaos_y:readdata -> mm_interconnect_1:pio_chaos_y_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_y_s1_address;               // mm_interconnect_1:pio_chaos_y_s1_address -> pio_chaos_y:address
	wire          mm_interconnect_1_pio_chaos_y_s1_write;                 // mm_interconnect_1:pio_chaos_y_s1_write -> pio_chaos_y:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_y_s1_writedata;             // mm_interconnect_1:pio_chaos_y_s1_writedata -> pio_chaos_y:writedata
	wire          mm_interconnect_1_pio_chaos_z_s1_chipselect;            // mm_interconnect_1:pio_chaos_z_s1_chipselect -> pio_chaos_z:chipselect
	wire   [31:0] mm_interconnect_1_pio_chaos_z_s1_readdata;              // pio_chaos_z:readdata -> mm_interconnect_1:pio_chaos_z_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_z_s1_address;               // mm_interconnect_1:pio_chaos_z_s1_address -> pio_chaos_z:address
	wire          mm_interconnect_1_pio_chaos_z_s1_write;                 // mm_interconnect_1:pio_chaos_z_s1_write -> pio_chaos_z:write_n
	wire   [31:0] mm_interconnect_1_pio_chaos_z_s1_writedata;             // mm_interconnect_1:pio_chaos_z_s1_writedata -> pio_chaos_z:writedata
	wire   [31:0] mm_interconnect_1_pio_chaos_temp_s1_readdata;           // pio_chaos_temp:readdata -> mm_interconnect_1:pio_chaos_temp_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_chaos_temp_s1_address;            // mm_interconnect_1:pio_chaos_temp_s1_address -> pio_chaos_temp:address
	wire   [31:0] hps_0_f2h_irq0_irq;                                     // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                     // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          log_generate_0_dout_valid;                              // LOG_Generate_0:dout_valid -> avalon_st_adapter:in_0_valid
	wire   [23:0] log_generate_0_dout_data;                               // LOG_Generate_0:dout_data -> avalon_st_adapter:in_0_data
	wire          log_generate_0_dout_ready;                              // avalon_st_adapter:in_0_ready -> LOG_Generate_0:dout_ready
	wire          log_generate_0_dout_startofpacket;                      // LOG_Generate_0:dout_sop -> avalon_st_adapter:in_0_startofpacket
	wire          log_generate_0_dout_endofpacket;                        // LOG_Generate_0:dout_eop -> avalon_st_adapter:in_0_endofpacket
	wire    [1:0] log_generate_0_dout_empty;                              // LOG_Generate_0:dout_empty -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                          // avalon_st_adapter:out_0_valid -> timing_adapter_0:in_valid
	wire   [23:0] avalon_st_adapter_out_0_data;                           // avalon_st_adapter:out_0_data -> timing_adapter_0:in_data
	wire          avalon_st_adapter_out_0_ready;                          // timing_adapter_0:in_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                  // avalon_st_adapter:out_0_startofpacket -> timing_adapter_0:in_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                    // avalon_st_adapter:out_0_endofpacket -> timing_adapter_0:in_endofpacket
	wire          rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [LOG_Generate_0:reset, alt_vip_itc_0:rst, alt_vip_mix_0:reset, alt_vip_tpg_0:reset, alt_vip_vfr_0:reset, avalon_st_adapter:in_rst_0_reset, mm_interconnect_1:alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset, timing_adapter_0:reset_n]
	wire          rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [alt_vip_vfr_0:master_reset, mm_interconnect_0:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire          rst_controller_002_reset_out_reset;                     // rst_controller_002:reset_out -> [mm_interconnect_1:pio_chaos_done_reset_reset_bridge_in_reset_reset, pio_chaos_done:reset_n, pio_chaos_reset:reset_n, pio_chaos_shift:reset_n, pio_chaos_step:reset_n, pio_chaos_temp:reset_n, pio_chaos_w:reset_n, pio_chaos_x:reset_n, pio_chaos_y:reset_n, pio_chaos_z:reset_n]
	wire          rst_controller_003_reset_out_reset;                     // rst_controller_003:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire          rst_controller_004_reset_out_reset;                     // rst_controller_004:reset_out -> mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	log_generator #(
		.BACK_COLOR        (26'b00000000000000000000000001),
		.FRONT_COLOR       (26'b00111111111111111111111111),
		.MIF_FILE_LOCATION ("./log.mif"),
		.LOG_WIDTH         (1024),
		.LOG_HEIGHT        (249)
	) log_generate_0 (
		.reset      (rst_controller_reset_out_reset),    //      reset.reset
		.clock      (pll_stream_outclk1_clk),            // clock_sink.clk
		.dout_ready (log_generate_0_dout_ready),         //       dout.ready
		.dout_valid (log_generate_0_dout_valid),         //           .valid
		.dout_data  (log_generate_0_dout_data),          //           .data
		.dout_sop   (log_generate_0_dout_startofpacket), //           .startofpacket
		.dout_eop   (log_generate_0_dout_endofpacket),   //           .endofpacket
		.dout_empty (log_generate_0_dout_empty)          //           .empty
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (640),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (639),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (10),
		.V_BACK_PORCH                  (33),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_stream_outclk1_clk),                    //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),            // is_clk_rst_reset.reset
		.is_data       (alt_vip_mix_0_dout_data),                   //              din.data
		.is_valid      (alt_vip_mix_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_mix_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_mix_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_mix_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	soc_system_alt_vip_mix_0 alt_vip_mix_0 (
		.clock                 (pll_stream_outclk1_clk),                              //   clock.clk
		.reset                 (rst_controller_reset_out_reset),                      //   reset.reset
		.din_0_ready           (alt_vip_tpg_0_dout_ready),                            //   din_0.ready
		.din_0_valid           (alt_vip_tpg_0_dout_valid),                            //        .valid
		.din_0_data            (alt_vip_tpg_0_dout_data),                             //        .data
		.din_0_startofpacket   (alt_vip_tpg_0_dout_startofpacket),                    //        .startofpacket
		.din_0_endofpacket     (alt_vip_tpg_0_dout_endofpacket),                      //        .endofpacket
		.din_1_ready           (timing_adapter_0_out_ready),                          //   din_1.ready
		.din_1_valid           (timing_adapter_0_out_valid),                          //        .valid
		.din_1_data            (timing_adapter_0_out_data),                           //        .data
		.din_1_startofpacket   (timing_adapter_0_out_startofpacket),                  //        .startofpacket
		.din_1_endofpacket     (timing_adapter_0_out_endofpacket),                    //        .endofpacket
		.din_2_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),         //   din_2.ready
		.din_2_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),         //        .valid
		.din_2_data            (alt_vip_vfr_0_avalon_streaming_source_data),          //        .data
		.din_2_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //        .startofpacket
		.din_2_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //        .endofpacket
		.dout_ready            (alt_vip_mix_0_dout_ready),                            //    dout.ready
		.dout_valid            (alt_vip_mix_0_dout_valid),                            //        .valid
		.dout_data             (alt_vip_mix_0_dout_data),                             //        .data
		.dout_startofpacket    (alt_vip_mix_0_dout_startofpacket),                    //        .startofpacket
		.dout_endofpacket      (alt_vip_mix_0_dout_endofpacket),                      //        .endofpacket
		.control_av_chipselect (mm_interconnect_1_alt_vip_mix_0_control_chipselect),  // control.chipselect
		.control_av_write      (mm_interconnect_1_alt_vip_mix_0_control_write),       //        .write
		.control_av_address    (mm_interconnect_1_alt_vip_mix_0_control_address),     //        .address
		.control_av_writedata  (mm_interconnect_1_alt_vip_mix_0_control_writedata),   //        .writedata
		.control_av_readdata   (mm_interconnect_1_alt_vip_mix_0_control_readdata)     //        .readdata
	);

	soc_system_alt_vip_tpg_0 alt_vip_tpg_0 (
		.clock              (pll_stream_outclk1_clk),           // clock.clk
		.reset              (rst_controller_reset_out_reset),   // reset.reset
		.dout_ready         (alt_vip_tpg_0_dout_ready),         //  dout.ready
		.dout_valid         (alt_vip_tpg_0_dout_valid),         //      .valid
		.dout_data          (alt_vip_tpg_0_dout_data),          //      .data
		.dout_startofpacket (alt_vip_tpg_0_dout_startofpacket), //      .startofpacket
		.dout_endofpacket   (alt_vip_tpg_0_dout_endofpacket)    //      .endofpacket
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (640),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (639),
		.RMASTER_BURST_TARGET           (64),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_0 (
		.clock                (pll_stream_outclk1_clk),                                 //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (pll_sdram_outclk1_clk),                                  //            clock_master.clk
		.master_reset         (rst_controller_001_reset_out_reset),                     //      clock_master_reset.reset
		.slave_address        (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                          //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                         //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                         //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                       //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                        //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                       //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                      //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                      //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                       //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                    //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                         //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                        //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                      //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                        //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                         //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                      //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),  //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),  //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),               //         h2f_reset.reset_n
		.h2f_axi_clk              (pll_sdram_outclk1_clk),                 //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),             //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),           //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),            //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),           //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),          //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),           //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),          //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),           //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),          //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),          //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),              //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),            //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),            //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),            //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),           //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),           //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),              //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),            //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),           //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),           //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),             //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),           //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),            //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),           //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),          //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),           //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),          //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),           //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),          //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),          //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),              //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),            //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),            //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),            //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),           //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),           //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),        //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),         //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),        //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),       //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),        //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),       //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),        //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),       //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),       //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),           //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),         //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),         //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),         //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),        //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),        //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),           //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),         //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),        //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),        //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),          //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),        //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),         //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),        //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),       //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),        //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),       //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),        //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),       //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),       //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),           //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),         //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),         //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),         //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),        //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),        //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                    //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                     //          f2h_irq1.irq
	);

	soc_system_pio_chaos_done pio_chaos_done (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_pio_chaos_done_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pio_chaos_done_s1_readdata), //                    .readdata
		.in_port  (pio_chaos_done_external_connection_export)     // external_connection.export
	);

	soc_system_pio_chaos_reset pio_chaos_reset (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_reset_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_reset_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_shift pio_chaos_shift (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_shift_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_shift_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_shift_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_shift_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_shift_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_shift_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_reset pio_chaos_step (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_step_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_step_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_step_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_step_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_step_s1_readdata),   //                    .readdata
		.out_port   (pio_chaos_step_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_temp pio_chaos_temp (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_1_pio_chaos_temp_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pio_chaos_temp_s1_readdata), //                    .readdata
		.in_port  (pio_chaos_temp_external_connection_export)     // external_connection.export
	);

	soc_system_pio_chaos_w pio_chaos_w (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_w_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_w_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_w pio_chaos_x (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_x_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_x_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_w pio_chaos_y (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_y_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_y_external_connection_export)       // external_connection.export
	);

	soc_system_pio_chaos_w pio_chaos_z (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_chaos_z_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_chaos_z_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_chaos_z_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_chaos_z_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_chaos_z_s1_readdata),   //                    .readdata
		.in_port    (pio_chaos_z_external_connection_export)       // external_connection.export
	);

	soc_system_pll_sdram pll_sdram (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~reset_reset_n),        //   reset.reset
		.outclk_0 (sdram_clk_clk),         // outclk0.clk
		.outclk_1 (pll_sdram_outclk1_clk), // outclk1.clk
		.locked   ()                       //  locked.export
	);

	soc_system_pll_stream pll_stream (
		.refclk   (clk_clk),                        //  refclk.clk
		.rst      (~reset_reset_n),                 //   reset.reset
		.outclk_0 (clock_bridge_148_5_out_clk_clk), // outclk0.clk
		.outclk_1 (pll_stream_outclk1_clk),         // outclk1.clk
		.locked   ()                                //  locked.export
	);

	soc_system_sdram sdram (
		.clk            (pll_sdram_outclk1_clk),                    //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	soc_system_timing_adapter_0 timing_adapter_0 (
		.clk               (pll_stream_outclk1_clk),                //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),       // reset.reset_n
		.in_data           (avalon_st_adapter_out_0_data),          //    in.data
		.in_valid          (avalon_st_adapter_out_0_valid),         //      .valid
		.in_ready          (avalon_st_adapter_out_0_ready),         //      .ready
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //      .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //      .endofpacket
		.out_data          (timing_adapter_0_out_data),             //   out.data
		.out_valid         (timing_adapter_0_out_valid),            //      .valid
		.out_ready         (timing_adapter_0_out_ready),            //      .ready
		.out_startofpacket (timing_adapter_0_out_startofpacket),    //      .startofpacket
		.out_endofpacket   (timing_adapter_0_out_endofpacket)       //      .endofpacket
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                 //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),               //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),               //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),              //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),               //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),              //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),               //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),              //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),              //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                  //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),               //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),               //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                  //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),               //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),               //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                 //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),               //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),               //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),              //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),               //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),              //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),               //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),              //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),              //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                  //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),               //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),               //                                                           .rready
		.pll_sdram_outclk1_clk                                            (pll_sdram_outclk1_clk),                     //                                          pll_sdram_outclk1.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),        //     alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),        // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                              (alt_vip_vfr_0_avalon_master_address),       //                                alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                          (alt_vip_vfr_0_avalon_master_waitrequest),   //                                                           .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                           (alt_vip_vfr_0_avalon_master_burstcount),    //                                                           .burstcount
		.alt_vip_vfr_0_avalon_master_read                                 (alt_vip_vfr_0_avalon_master_read),          //                                                           .read
		.alt_vip_vfr_0_avalon_master_readdata                             (alt_vip_vfr_0_avalon_master_readdata),      //                                                           .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                        (alt_vip_vfr_0_avalon_master_readdatavalid), //                                                           .readdatavalid
		.sdram_s1_address                                                 (mm_interconnect_0_sdram_s1_address),        //                                                   sdram_s1.address
		.sdram_s1_write                                                   (mm_interconnect_0_sdram_s1_write),          //                                                           .write
		.sdram_s1_read                                                    (mm_interconnect_0_sdram_s1_read),           //                                                           .read
		.sdram_s1_readdata                                                (mm_interconnect_0_sdram_s1_readdata),       //                                                           .readdata
		.sdram_s1_writedata                                               (mm_interconnect_0_sdram_s1_writedata),      //                                                           .writedata
		.sdram_s1_byteenable                                              (mm_interconnect_0_sdram_s1_byteenable),     //                                                           .byteenable
		.sdram_s1_readdatavalid                                           (mm_interconnect_0_sdram_s1_readdatavalid),  //                                                           .readdatavalid
		.sdram_s1_waitrequest                                             (mm_interconnect_0_sdram_s1_waitrequest),    //                                                           .waitrequest
		.sdram_s1_chipselect                                              (mm_interconnect_0_sdram_s1_chipselect)      //                                                           .chipselect
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                           //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                         //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                          //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                         //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                        //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                         //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                        //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                         //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                        //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                        //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                            //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                          //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                          //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                          //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                         //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                         //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                            //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                          //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                         //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                         //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                           //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                         //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                          //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                         //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                        //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                         //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                        //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                         //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                        //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                        //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                            //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                          //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                          //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                          //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                         //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                         //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                //                                                     clk_0_clk.clk
		.pll_stream_outclk1_clk                                              (pll_stream_outclk1_clk),                                 //                                            pll_stream_outclk1.clk
		.alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                         //         alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                     // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.pio_chaos_done_reset_reset_bridge_in_reset_reset                    (rst_controller_002_reset_out_reset),                     //                    pio_chaos_done_reset_reset_bridge_in_reset.reset
		.alt_vip_mix_0_control_address                                       (mm_interconnect_1_alt_vip_mix_0_control_address),        //                                         alt_vip_mix_0_control.address
		.alt_vip_mix_0_control_write                                         (mm_interconnect_1_alt_vip_mix_0_control_write),          //                                                              .write
		.alt_vip_mix_0_control_readdata                                      (mm_interconnect_1_alt_vip_mix_0_control_readdata),       //                                                              .readdata
		.alt_vip_mix_0_control_writedata                                     (mm_interconnect_1_alt_vip_mix_0_control_writedata),      //                                                              .writedata
		.alt_vip_mix_0_control_chipselect                                    (mm_interconnect_1_alt_vip_mix_0_control_chipselect),     //                                                              .chipselect
		.alt_vip_vfr_0_avalon_slave_address                                  (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_address),   //                                    alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                                    (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_write),     //                                                              .write
		.alt_vip_vfr_0_avalon_slave_read                                     (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_read),      //                                                              .read
		.alt_vip_vfr_0_avalon_slave_readdata                                 (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_readdata),  //                                                              .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                                (mm_interconnect_1_alt_vip_vfr_0_avalon_slave_writedata), //                                                              .writedata
		.pio_chaos_done_s1_address                                           (mm_interconnect_1_pio_chaos_done_s1_address),            //                                             pio_chaos_done_s1.address
		.pio_chaos_done_s1_readdata                                          (mm_interconnect_1_pio_chaos_done_s1_readdata),           //                                                              .readdata
		.pio_chaos_reset_s1_address                                          (mm_interconnect_1_pio_chaos_reset_s1_address),           //                                            pio_chaos_reset_s1.address
		.pio_chaos_reset_s1_write                                            (mm_interconnect_1_pio_chaos_reset_s1_write),             //                                                              .write
		.pio_chaos_reset_s1_readdata                                         (mm_interconnect_1_pio_chaos_reset_s1_readdata),          //                                                              .readdata
		.pio_chaos_reset_s1_writedata                                        (mm_interconnect_1_pio_chaos_reset_s1_writedata),         //                                                              .writedata
		.pio_chaos_reset_s1_chipselect                                       (mm_interconnect_1_pio_chaos_reset_s1_chipselect),        //                                                              .chipselect
		.pio_chaos_shift_s1_address                                          (mm_interconnect_1_pio_chaos_shift_s1_address),           //                                            pio_chaos_shift_s1.address
		.pio_chaos_shift_s1_write                                            (mm_interconnect_1_pio_chaos_shift_s1_write),             //                                                              .write
		.pio_chaos_shift_s1_readdata                                         (mm_interconnect_1_pio_chaos_shift_s1_readdata),          //                                                              .readdata
		.pio_chaos_shift_s1_writedata                                        (mm_interconnect_1_pio_chaos_shift_s1_writedata),         //                                                              .writedata
		.pio_chaos_shift_s1_chipselect                                       (mm_interconnect_1_pio_chaos_shift_s1_chipselect),        //                                                              .chipselect
		.pio_chaos_step_s1_address                                           (mm_interconnect_1_pio_chaos_step_s1_address),            //                                             pio_chaos_step_s1.address
		.pio_chaos_step_s1_write                                             (mm_interconnect_1_pio_chaos_step_s1_write),              //                                                              .write
		.pio_chaos_step_s1_readdata                                          (mm_interconnect_1_pio_chaos_step_s1_readdata),           //                                                              .readdata
		.pio_chaos_step_s1_writedata                                         (mm_interconnect_1_pio_chaos_step_s1_writedata),          //                                                              .writedata
		.pio_chaos_step_s1_chipselect                                        (mm_interconnect_1_pio_chaos_step_s1_chipselect),         //                                                              .chipselect
		.pio_chaos_temp_s1_address                                           (mm_interconnect_1_pio_chaos_temp_s1_address),            //                                             pio_chaos_temp_s1.address
		.pio_chaos_temp_s1_readdata                                          (mm_interconnect_1_pio_chaos_temp_s1_readdata),           //                                                              .readdata
		.pio_chaos_w_s1_address                                              (mm_interconnect_1_pio_chaos_w_s1_address),               //                                                pio_chaos_w_s1.address
		.pio_chaos_w_s1_write                                                (mm_interconnect_1_pio_chaos_w_s1_write),                 //                                                              .write
		.pio_chaos_w_s1_readdata                                             (mm_interconnect_1_pio_chaos_w_s1_readdata),              //                                                              .readdata
		.pio_chaos_w_s1_writedata                                            (mm_interconnect_1_pio_chaos_w_s1_writedata),             //                                                              .writedata
		.pio_chaos_w_s1_chipselect                                           (mm_interconnect_1_pio_chaos_w_s1_chipselect),            //                                                              .chipselect
		.pio_chaos_x_s1_address                                              (mm_interconnect_1_pio_chaos_x_s1_address),               //                                                pio_chaos_x_s1.address
		.pio_chaos_x_s1_write                                                (mm_interconnect_1_pio_chaos_x_s1_write),                 //                                                              .write
		.pio_chaos_x_s1_readdata                                             (mm_interconnect_1_pio_chaos_x_s1_readdata),              //                                                              .readdata
		.pio_chaos_x_s1_writedata                                            (mm_interconnect_1_pio_chaos_x_s1_writedata),             //                                                              .writedata
		.pio_chaos_x_s1_chipselect                                           (mm_interconnect_1_pio_chaos_x_s1_chipselect),            //                                                              .chipselect
		.pio_chaos_y_s1_address                                              (mm_interconnect_1_pio_chaos_y_s1_address),               //                                                pio_chaos_y_s1.address
		.pio_chaos_y_s1_write                                                (mm_interconnect_1_pio_chaos_y_s1_write),                 //                                                              .write
		.pio_chaos_y_s1_readdata                                             (mm_interconnect_1_pio_chaos_y_s1_readdata),              //                                                              .readdata
		.pio_chaos_y_s1_writedata                                            (mm_interconnect_1_pio_chaos_y_s1_writedata),             //                                                              .writedata
		.pio_chaos_y_s1_chipselect                                           (mm_interconnect_1_pio_chaos_y_s1_chipselect),            //                                                              .chipselect
		.pio_chaos_z_s1_address                                              (mm_interconnect_1_pio_chaos_z_s1_address),               //                                                pio_chaos_z_s1.address
		.pio_chaos_z_s1_write                                                (mm_interconnect_1_pio_chaos_z_s1_write),                 //                                                              .write
		.pio_chaos_z_s1_readdata                                             (mm_interconnect_1_pio_chaos_z_s1_readdata),              //                                                              .readdata
		.pio_chaos_z_s1_writedata                                            (mm_interconnect_1_pio_chaos_z_s1_writedata),             //                                                              .writedata
		.pio_chaos_z_s1_chipselect                                           (mm_interconnect_1_pio_chaos_z_s1_chipselect)             //                                                              .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_stream_outclk1_clk),                // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (log_generate_0_dout_data),              //     in_0.data
		.in_0_valid          (log_generate_0_dout_valid),             //         .valid
		.in_0_ready          (log_generate_0_dout_ready),             //         .ready
		.in_0_startofpacket  (log_generate_0_dout_startofpacket),     //         .startofpacket
		.in_0_endofpacket    (log_generate_0_dout_endofpacket),       //         .endofpacket
		.in_0_empty          (log_generate_0_dout_empty),             //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_stream_outclk1_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_sdram_outclk1_clk),              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (pll_sdram_outclk1_clk),              //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
