��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW��3��+�M|�Qb"+��#�g?	t<�	��M/<��eg;���B�`}Mh�0^F
1��<%��a6�t?�n�+�hX�o>�AJkG�iQI���*@)������f��%��Ǟ�H� �a�C��|�� �P�Y�v��K��b��g�?��w� 1)��9Қ9��}I,�/{����OF#(�����\x�XCמ'�è+C��4L�6
�e6�"�}�y�!�e��)��ܨ0�E;��]Q�rqR9ڥß� �#�	\V��& #���������h0���cx7I�%�a�(��n3�8~�Y�@��Qg[��Wl���5nRo�ȊF�I1�n؂����ި�+"$�ߏ��?%î���a��o����XN勞����1;d���>p�	^:ƿ��	�1��\R�d���(�"pW�A��6��6_)_!���_x3�I����$���q��^�퍨av�������+�\�P)�'c�bt>3b@T{�����
��P��B%�S=X)2�_E����_SI���͢z�:ұ�����d�mu ���u�[`,� �Z[gw��LoI�������$"nogg�W��P.��a���:4��`��,Џ}�_)!����`mK�rg��nD�����^��vT�-]$�u<��N��+���9�)��L8�p:��O�oO>�J�~M�*���M��P�*?���#�"�I<�
9cW�}��m��bu�ja�Pu|����ΧM�-����&�3�`Z�΂꺾��V��H�&3���ܰQ���
�g�LĴ�,�C�M�:���JQ�Ϋ��u���8[J%"��b]���?uj�3C�.��m[���!���b�:t� ��t���X8T�eF�5��Sє�!@�f�|�bת4�U�>܏>����9IWP�(�~0Gs�`͏8*�3�ɖ�/�t�$Od��ϱ�� ���7:��	��"|3"���L�������ǅ+E�N� /��APP�Zؓj�S>v�5���Xŝ�`�U�	K� /u�7hЀf��cj��/h�����p��F1�3rF�t�^ϰ:]����3�q�:��������Ԑg�$�����!;��+�L�Bp�G�9׵�C/$)�ftq�������}O7�fq�[El�[R��;Hf���
xM�G﬍�Q�E��i�N�ң��v�G�&��QꝔ,�*���Az�w
/L��d(�?׆2:���kh!.���Y�Z%oQ��ddD��!��ªذ��o�����	�B	i+��57�3C�t �rx㡶#IR�[=�Wg�������IMex��)W�6���;���u�?��N��xmo�H�c&_y�[�Å��<<
�0`r�ߤ0������p@����၍ ��'JZ�r�v�j�����!X˓_"�i$�^_\b�im;P�uj�*;����g�'�yT�h6!�.�A:�Rk�˝��h"R�޺�	���?�5AoM�⣨�$��c�7�N1 ����Rc�4�MH�o>�=�YQ�(���d ]I��w+�CK��v-l���c��<���nWBŻ�'	n���t�Z2j`k^���7j����J{$ �}��Y�*��{�e�%����g}@V_���z]��R���q0��DD���i&��g�K�/�E��]bO@�>�ޒa���>��ŧ��	y�=&8MJ�������ڌ�~�Y�g)���k�wsŮ���uh��i&�?(��'���Iυ�F�;	,v�q�
G��8�E<}#%�v�\j�^g޹�7b�� X��C�ߥ�!n��q�K���Y�ɸtv� �?�"ίk�N�M4��V�"&AJ�`
�!.������E4��T}pz��w��T#N�ܕ�x���<j	�&*)��]�V�C��K�f�V���WIt.z�|�$��-H�\U�e�(WY�}�ñ�n�7�փ��c�����3g8�`��]��2Ӭ��p|l���+A�+|-y�R2��J����q.$R�~A��$��.g8ݕ���Uy�TG��ٕp��ȷD�)�?�����+/m�KI!�O��*Yn�y(�}�fF�V�n��Z��pǚ��7Vl ���x�T�M$� �������ڢ;#
Ba��*�>TLSI����:Y[���t�VNRB/W�M�Z����y�;��'"G���/���y�=`�U��|�p�*ޏ]H���-��w>W�`Gj�AW!��&C]~>��x�]
N��3�������מ*�_(ƃϠb���#������y��@=�=ʣX�{8$"����GD�Zai�RcԨǤ��9d�Q�%Il�T�E�- O�o:a����?�d�y��۝��&�RQ�uS:֎�(�2�u�a�w�k� y^�k�<Y�ͣ S�y��6��k!j_F�K�~���c��@Ѷ�Sr�ϴ��mZ�#�������"�,)Q�u�<�.N/쯁0��S�>�5!�V'�M0��j�t7+6�+~��N̺lѼ�K�[s��sb����K��>�ZS��a����	��]�32n��N�%���I�E�b4��:V�|F��f��+���{px�tK�i���%ܑ� F�V�1TW��.9�puF{vޤ{$0�M�(s�� ��El��L:<w	�2R�VJ���}���9�q��SJ����QR, �lom]�BO&Ҏk[Z��4��-��:��t�C_��k�f)�G�U�!�+��V�3�]:��$�o*�ڠ���
��p�Xe�j+����hc���%h����v޶�e��G(��3�ũ�n�s����`&�7;��ee�N��7��M��Վ���C��q�����	��/�zU�_�<�\�p@����I�J�M�)f�%P��wd~�=����8��Ai(��oj� oHw?Fu�4�ƫd�g�L��[��Jv쵊�����M<&��6`�`�rFi�8�'����`���*�(ϖ�5L��Ŕ��� z)�qŔ���u؟iQR�x�� -,�!0T�m5{y��\���{R^�g�n��n6�z|yc��6�  £[��R 7t�RcL~�<�,�Qz������Iq7�����N���fG�/9T��Q��k߻:_N����1'�}��6�A��,=�p}�#�5�b^Ei����n�bFVR�|��K���N*F� hxLAI!W�m=�RM�H�70�B��m�����N)�_!�1��J`�8��b7L��%Ъ=�*���3i����bSi�f@n�Wx�Z����q}�?�!��ϙ9-�Rׯzr�c1"� w̜�J�D^|(9f�q(��A6��V�����Ē����_�)R��[�hDGhռ[6 ���*�3W� ՗�$�X�m����{��������$��9�ӄ�:����Ed��{P3��/�j�X�\^�Am�9���wϬ�n��I�Ѝ�bf�L�H��,�9�� ��	7Xf�_�a��W���x�uS�[�:��x�嗐/��%�+�/T0�������9�-�2��K�g����z7*����T��7�aI�AҢX�%�e��w���n�uV�������@(�ޑu�����.6԰�6����Wʏ�3@��7ؕ �j�2���M��$�<Ec�~O�e{���8JJFw��)�� szfL����+N�#�Mk�� ���1�f���� OX	��;�UI��Z�2�~�ӀF�
n��	�nE���q�7ؕQ���kb/D��A��9-�&�g���9�4�ݎ��zS��?x���}�\��o(iu���u����C���\���R�u(�D��"�	��#5�����~�Z4[D*�A�H�
�ņ�E�{�>�hV�����l���mɚ�GL{r-d��q��� ��Uf3ַi��7E�v�S�;��b�욺{_e?I`���%��&i �l�jKtju����b���=��W�K��'�yJv7���"2蚰P�,�-L-�	��u��!�����b����
�N�c^��%3�ķ|����C���@��Q/��?�4}ǽRNj%V����pa8��|z��$8ݩ���գ/s�UǬ�Db7���99��:�8�)�Vm���4��^r� J��A��b�i��8I��4{]����|�zZ�	���ׅ���!Ox30F�+�C1�-�����֏�{����<S
?�4�%u���G�����Eb�aL#�8���.8v3�f��S�I'ꫠ��G�n���xmLġ-8�ٗ�]��:=ܽ����{���J�[��ò� �m�������uX�(���hu��v���t�_��!B��%<��Zn�ף�4v�.�	A�Dr� ũ��~���N�n��Ӣρ{���DYM�_T��U��U��K�5�e��7j]y�0*�*��9�pҲ�T�T�����_x.���<�T�UZ��D%l=`]�Nc���p�]Ղ�n��q�5׃/]�W����5�[�ڲ���\e"��U~Ȕ�:��v}sqk���DqPm�bn���Lys�����p��l�?镡���C�^�)�(Ƅ��Er�@�;u��Q"a�\#oa�/>X�fISV٢7��ԁN{E�lCx�a��I` ���y$�.����� �|��[`D�m�#�/�Q�ٱ/�� c����ײ>4�o%�ӽz8���	Ob�0�nxlf5���G�A�h�&G]sE�'u���Pg���?��E^���$��-�����'��)`tɞ=?A�I�Ck�7>a�1s�dĮ�p�u��J�eJب8?�^S�9���]չ��ʸ�����~�$U�"m�}~}vb��6��Ak��$c����*�K3z=YxOQ�E���8����۹>T�DaJЈ� a�� Z�4���+����a�e��zr�x\���Rk)-�3ϣ�1���5�{�GBڃ���2^EĔ�4��%�+d�!مtA�W*G��t��sUJ��'�.�<�X�`��~V�.q�#?>sxI������<kNtg�/+�ح~���N��6��B��hI�$^z�'���cA �Hy<�
.��{���e��&�q��8��Z���#h��z���4s� 2-�!��M�M刭����
�=%�
+]b�H�](�r�q�Q�d9�N�¢3ْ��r�5?v<#���t쎷�EH�ցlf~3_o��Kc5�)��RuY~�ң�EqҼ�A0T�i������t�v2�|J<����R�W�%v�V/<��qmu]��c�M�%7K��>��⧩(�X���:N"���L��Kcu_1"���!��Nq���N�b��j��p] ��ʊTl����R����!���5 �=���Z��NA��B���I�;��CE$��N��0{��!�l���u9����\`Z����6�>V�hV*��������'J�ۄ�{T�EU\�A����*����-؄D�� ��ͦd�E��/��ɮ�/�/�N�֕<<�}\yC'g��1RE��;3�f>N�Gr���Vlc.�RĖ3c�u�f�Ȓ�tO���.+�*��҈�_��i�eu�q�b0�~[<I�BcՖ�4��.AF y��g��VK�Qi���z׳UJ����9cz��ΞP� �SP���x�L�i������WoN[��-.� F"ƌ�#M�A��B���5Vq�J��*虘��UZ�E*t��3�v�qRv�P��X;BKK�s|���%Qf|/�;�C+X ������E�w.��M�X�TaR}���}�)
���*-���b	�$�^7{�͎m�
l����2Rx�%�R&�	��8�0�ў�C���jq�3�d��,��g��_#(��@R;k�O�~VgJ��|��ޱ�GYp���,غ���n��Y}���G����M꧶%;	� n�U���ӵs�ڇ���&�U� �e�s�/�x?v%>#��#��u�L6_�z��[��+R2���oE�ց-��8:-�X�%����&��M���I�nSԤ��gT<�)���������=F'���SM�k�J߯��aN�*�ɺ辗~�`=��X��;�/�D]`so-$�L!�g���b5��Q���k�:�PM�0����d�'N��T�m(�A���C7�_��#t-��Ұ9��,9Fs�CAi���ޫNi)����a����(E/�&�5��3(O4����2��M��&�2V�\)�nE��S��<9�&�
z��DW���:�l��R�Y��
�%VsC�x�Z�X\�Ц�O^F����ŭ���"-؀ϙDǢc�m�����@��#e�$s�<��]��G�ܰ���u �]6iK&�V�t_��=5��ӰV�ZG�m�
8F��J�Hed0vr�	}�o=TL�d�C��{E�$M�e��J��XmZ� ��)\.�ܝ��UdR�Z��B���=�Ǝ�|�����[tDe���7��`i_����6��R/�Eoo�*XN돛y\ځ����M�R.�e�%��{�ǐ�ٞ̑]���� .D���J+r�M+��w��ؿ�A��C(���DXT�&�k9	]Bs#�?M&� �:��_�e_HLLR����4Y���t ��P��x>k��R'"�rɸL�H��ߑ��U��DCc����h<zq�g��㧬��B~��q�~
>�`d�#c��uIL�� �s���� ��X�O"�ྌ����)	�QP����2���3d��\���~u�J��+�㧛z�w��N����G����kއ������̲c#VZ�.2D��t���	�D�Rݦ�t*Q�O[�g>�㰠��\v�,L��O��1^��l���>m��;WM����H�� m�wS�+Q�K�"��֜����u`SY<����(/sܮ�Kg�*e��؃�j��b�E�5"����\'s�7D��:e(�Jh�z��o�@٬kdR-}��R؝������z�v˹W����wm1�Q��(/�|J����α97+D����鵛X�����`�Ҵ��Zi)�gs]��_�"Bdh����(�ѡeL��e�-���7�/'�y���Ή� ʆ��FBy,dѶV���gŏR|�R�;���ߩ��|����M��C�E3�h�`�h���z RGtP��s^蚑"�����kw�%�[W>�^�J�ff-��������
�	+q\���PǵA�Z�d9�T��2�<�����u�mה]UjJ\'$<x8;2Z)h��4Y]���-�1�`u��qr� ��9�_Hv�08�r����"��MY}�J���	���U��S\-��
��m�on�������s��yܻV
�+Y�r��-�1�������Q���i�! ���v�	��_?�����E���uvN��?z������/>ã�<�Ì�uI�!�{��Pޭ�� �z�>8�� � �<Q�Wf�_w�B������q�d�i����O4} ���u��� ���y��]�����f�RU�G�������5�K��!�je�8�/*(wv�_x��&gx�����<�7n!���#��^��Z��*"�dM>���p�5E��e�n�ϟ��yP�r]�%��+ ����JNF��b6���������U��J耛{]d���\oU��5��,c��7n�삧�⑻^����^K�����%jS�?r��K)@wtL0fKhly?t�<�b�o�c�[>�V�c��&��b�]�ѵ�0k�K��6�Y9��A"+�{�zɩM"�Q�*`Y��K�o�y:�	���d�I� j� 멩q��ʝ��ٟP{�!���H)��1�E�SB|ә>*��q��rj��~d��#}w����T��8�������� �u�-�RV��;�������1(S��]w�Ǥ�n���3��K�����*��oV�+ܟ��h[m ��S�}u�ę����H�#3�8G@Ä1B%{�U�&ZO�x��h�!�WG|�dռ�r���e��I�DL��\����>��������Myx��M�h���4�a6�E��ܞ�lEh^���Zy9<�/P�p�B�a�hfϘ�^�o�/�=B<<��v����I�������0?T;[�g\�k���Lh�Yg�����������Ӷ�ன�}�����W`�#�����0L�����[� ��|�e�����>��M�_�~|!`��G뇁�A�>�d��/VjZV��I\թ�&�R^�L��w�kI�x�X�\�xoPR
>�Y�j�H�gPl����XP �{-��S�!(o��}S�r��azDD�Qr� J\h��m��°-��3�zn��䣖�M}�K�:,��>�g�1�B��7�t��{��FHI�;�{³����Ň��/�(�,��J�g�>�ϲq��¹fKY�%8Ċ�7��F�|�Q**B���㯨O%�{����R���c���:2�M�N����w������$<%�,�.�N��@�`� �pp\a�&2'�Q~^
+Ң�e�u�?�t<0�4��#�C�������:��(��Nm�1��m��iY�w�J^~�2��C�5�����N0!��yY'l�G�A��Ǣ�^!(P���<(�>Q��e'gp���3��#S�=n�h���ng}�<iYYU�A-�E9�0��'�|�> ���P�o�]��!�I��}ě���z,��ڷ8�'�� �k^s1��]p٭)��9�?cm�dv��\xzq��Cb% �*)���K������>����븭�b�����;`�<m���G���ߨ���D%���p��(l�X����3v��-�gN�'�O�ػ���:n%��cf*C8��4\�~ҖC{Ř��).�Q�x=/hz�jc+{�X6�e(〜9H��c�;���ah8�^�(���(6���&��&����$�� �BRU��N����ۄЩ~97 ��O�ƴ�o�q�艹�Hci����8�:d�8���͜��U{>���p��@��f��y�n$Q��4[
���V�R����6Qi�\���yF�ۺ_��2�G���6�˽�Y�w(JY4ʩ��g�7��]L�4�}FBpt��o�[^�I�d�|F���sX*��m��[�-��_����_D��^tUTp�98�|F{���ƂSc����u���V����#3؞t��	��p1�R�7��U���d�rdԎ��T9@�_�mQ��A�v�<���v"�K@u�����q������mX���>��X!4�VqE+�}��ã��Z6�n˰���a��85��p,�m ь�H��Q �Q͌��.D�Hg�̵�k����/��}���m���G(zd9G<V���J���r�aF凘h{H۸a��������^�d�9��U"ר7G�Ũ_�`R�<�　T���؜����?RBb2�ʯz;��~�Ş;D�Y�A��+v�ja��@�𲫓�ANԅE+�=�i�.�V�m1J�p>�O4���[˜�����N;`��;��]?��*Kww�~�'-��k1=�]��FX���&*v�X����PjD���TZE�Rn�~�)�jzQ_%�m�G�0Ej�Zl��2y��d��H�)��&̵0`�+E�tHД�#+���>���wk>�F�T�稕��x��]=���v!��0�֌�v��i(����ڄ:Q�{�T����6F�c��"ύ8�P/�6M
HR�A^��`�ԭ�+�^�^��DGÜ��mƐ�N� �e�z@��ȅ��]���s\D�<B.�n�N7I�����@�& ��j���gD��l�I�@�aO�ǆ5z��	�s��N�*�nq�G��)dx�ܲ�n�̘T�� ����wՀSW���{G\]�i ����S&���Y-�n��G6h���'߹�s�����*�-��s\{���7$'ݲH��H�x�nG!C�Ŏ}��������F�Wf39
��*;Ҝ<�iwm2\�5�q-�?���y��!����1���Zvs�� fV���/�{����LC��aBQ�� '$'Z��[���\&ՠ	�"(�J��S�/����Z�~l��C縣	,��C���ׄ��n�`�����M�B]̷}Ǔ�xR���ꤑ.����m�v,�%��<��-ѸI�dky)G� ���g�V��G�).By��M�YP� �z�c��v: ��o ݿG/��0v	L-7V��{{0���/e��<�:L�8VTđ�-8��QH2|�~��p
{��P���`v�����̳�k�������@�xT���|��I` �/Z�AFBQ�X���3kk�T�Yt����ň'�N�-)F�s�����6�w	����:m�b�;��Ԣ�*�:�i*eD���6��4�2������֏�C	f��_�ۣ1���Q�N�b�#r�N-|�Lu�i���O%�N3��6Y�c��д��TE��~g>�᫩�������J����'��0&��9�9��%���ӤQ7�*L����":F�棆q��B�9�U�*hc�X��Pm�����T5|��3����z�ФT+��>v�RUJ%����R9Ń�J�^��zAV[� b6.}�]�a���
���,s7D����s�Ȣ�\H1ԩZ�px_���rV�I���β�X0hM�A�էȘ�։�ˈ�/��7�v��0�'���!S��Vb���s�_`>*#@�|?T��O��¾>U�&����X�(�VQ��X��2Z���1�$���5z��8��H��`mQ�g�##=�彡-7+�=�ώ��]7���b�zO�*<u���Խ��®�զ_x��&����hl\�1����"K����^!�Hd�DGأ�y{�QE&B�KC��������qp����"�W?�p���V@G�����.�'׸��0��}n�zr��'�/U�/��̶ӆ��x-�ۯ��ArBZN黩���Ϙ9T�4��k�w�,ȋ� �}��@P��%�:H��kp�3p��{��ĭ�\���]@%Yb������+�g nCR/�v��ߚ�v\�w5",Ov
�A��V���a{����G��vw����5���F��`�����15�D�_�G��N))qѤA�0��8�,�������+d��h�������Y�����*�sj	>0w;(�1�r��k���~�;�GL4���jb֜��cw�wD6	I�3��H�s���NiX�%�o*� �12B��'Lt--�aNs^�@���KC�2���S fKE�/��U��zG����aZ�w^s�`!�"��*�L���C����;=?�aQy-IN��K�I�(�e�v} r�Qm4�Q��aˬ��1Zb��
�)@7y��4t3*��ȳ�lY�?�</c{��	��M�#]�b�G�A!���g�@�
�m��i�jF��`�q�iS��~��9����Ox&���l�����/��U�q[+�P�)P]�W5V���Y�
�L�}���Ɲ��f
��!At�ݝg3&<O�ɻ�DƷ�z�[cOu��- wUjI����!��'Q�*H���F������\�}�����W�5��kIS��=�����K��1��˃�jh��񺫯k���2ᑨ���,���Js7WL0/�����AďT�܇��X�>w� �xv���s�.z'�g؟>E�b�V��e��D�V�<F�&�F�d��N���&�bQ:2-��oR��J����I��G��x��x8`=�&yX�A��D@���f�	
���m
�VJ��Fj��x�$HNu�Ne��M�F6뽊3����:��&��̀�5��(�-��L�:�s���7+��		��� W�%d)\0������b|�癚웕�0�]u�"���W�����I�� �|���Yi����zE! ��w�x��j���S10UNb��Rw��aL��V��Ѕ5
Ns�����P��Y`���@����+�2q�/�t��.o�J:O|[���iF�T�]�yI�$A&(�2/�Ħ�-&A?��I�8�fq��Z���X����#���{�H�{��݇7��#R���'�n�< QeJ�t�<܄B=��y�R�Y�ؑg|3�����10�����Ϟ/!3ڀ��K;��T��m�a��N�.���I�pt���!�A�o���V�po���A�_�g��E��z����@ޑĞ5b��YO��mTH60�ؔ�D�����	uF�O$�a��)�;�YH���RC�!�踜��� ��B���tJG��Ft�&n*~�F�}g�5�#?�d~��
u{V����,~A������3BT%%��1]��u����h)���?�g���O�Q|s�N��}%�6��'���:`����bu�)�	_�ȅy�Ķa	C�l��c�a+F}©
%�3�n_SǼ�~�d���|/Kߵ-_�	�]�L�|#���e�ɩ�vnU6��W���P����b���l6�0⌋:W�q���9��4��U\!�>d���H�S�~���´����x���A
F.>��kV�2�y�/l�:�l�a��䤡ȷD�EtE�d$�,���/q�G��O�<��!Lg-�
B0���94M�����MG�6��Nh�.��'1��.�Is�����o��kT;�F ��CV�:�	nIr�Q��v�/w�`�M��A3��D��ʣ�������c$Wb�=�h̋�����B���;L�<�4������H�T�K�D��ӧ1��|QGf@�K	��H�_I~ѤrD�S��)��̟����%A�Ȗ8�AjS�v��s�I��5��}HKC�&�в�E�x7�35��-²C���<P>�x�1�2�~�6�)�?p��mC�7�S:=P�ս���o|b�=���9$�C����X(��N��E-Z89 5����x�O�*�>旕+u�-�;	�vWT'����B)		��b�U)�:D� &bX�P�eR˵k${�{�X6ӒcS��}�*R�㮥܉�A8�����BxQ⥞�hy�ý�׻D�-�}��al�/�d�$��"�E���8@g��gSn�9�eC�@-O�� )že��S�<���>*�T�����@�9�������H٨�u<5�V�"�>�����͎����-����M���J���w���:���W'/�h/�G�!�u�t�Q����3�Ym��m������$3������+�N9��Hi�m-��8d1���Y��3Q]H�	����a�A�e�^eKَ과7��V� �)����ȿ��K�H��|��3�-1�b����Ⱥ$p<w���p"������D���zM��ש�O:��̆wy��_�E�����_��e���wP3��L�)W@��d�	��e�?�8жB�I�����_~/B�Y;_lڋ��h
�����_Ƭ���M�-:H'����e��t������������'�ϧ>;$Ýɳ��[�e�����r��	��84�B��������v���d�L˒h�bYV�'��Mqu�i���<z� m�oa6�N^�ŭ�h��{��2�#���a@έ
IV��'9��`�L�ïsc\�����-�V��ǊE�$c���P���8mw�;�o{̃豋��c	S�V_��F�[�w���V]��ݞ��sv��)�Q�*R��w��VQ���':ǯi�Ļ�F�#�4ϻP�N&)f0�)���,2J(V��^�mox�en8^(9��N*�1'O���/�RDωR�p���E�R�O�N]�'V�i̞q�<��]	��O�apV!Z �y�sQL������:��F�M���_�_��W
��e�+����i��C�2�9����&��A����`�e�1�~���v'�eo;��U�Ί�D�'Uz�|m��� ��<���ޟ�[ �����7�|Fz(����|&i]t�����EY;	RD���	��'S"ƭd�Q�"Qᚣg�����[���
y�Co[�9�jT�� b.g���(5�G��M�(p/$���K��`�oi�����s7PS.l-�cճH�#�2�-a���|{���h�l<F������S]Kp�2M����I/sQ'9����S*��H��ύ�G��-���#+� �QxW,,�H٠��5|�ܧEf[�1pt�(?�-_:i��d4��y�8��e�&G��)f���O�v���̖�N�+�T�r��*�T���r�[��l��!�:B2�l���v��Mhq=�,tC���F?��Ϳ3%�/F��SP���O&;�,���/�^?�Р�i6aКp�2_S	Ğ�8$-���L"V���P���z�~�tlU%Ļ�1E\�Xj&�fWـ�I�x�.���ѩ!7FOd܉Y
�R2�n����������ܤS���&.n�.o钳�E#G��g5�u��C�����qR���N7�iV0�of�C�)v���V��[!�:0���r�kɫ�A��,-v�un�So4+]��-߁�c6rͺ�7�����H+��Ӫ��O�c��ņe�P¦��f���D��]C����ګ����sv&*J�H;��?gk?V�2#à�
vD>�S��i`� vz4a����wc#���k�������S0([7����x�܂�x`�͟k=�ٓ�<��b��d����i���GI����#b�����p��`�Y�ņS���Ίu�p0��h��|��V=�שׂ��OU�Rd��sR5n��TVN��w-�J:��@����)���$S��r�a�[���ƒ|���V9~E�%��z��\�Z�BŮ0kT"*�d��@!B�����*;��L6E^4�eIտ6*)//�uy�&F�x��(I�����2��
���Dl0^Aj��ɔ� �W� �ޭE�lfA��n�|.L 72	�uc��ߍ��(ܦ�d�?�<�w��`��4nt��k��mm,�B��69���b��4�sA�mc̣��~�e<CC��~2���p�L��[�ƪm,x�[�w�Q.����e�wyW�H�O�x�DԲA�iJP=$&���D+�(/��t:.��L��T�`g�JJV6��r�H�����X\��v@�f,qЊ&�^ ��Rki��
s&x��u��v�q�Z�B%�	8j�%���POY�P����4-���R[i�/�2pP^()Y�$AT��5I�h&����];�GQ�T:��ױ��F�/z"cZC��`����^��JL	l�^�a�ʟ��am���v�����+
�g;y3oN���7 ����ZA�o��K�C0ͬ*ѩ��߇8��|]����m�4�5�,&a#������ki�C�ب��w<[pD`�v��>�]��w�u����w����cn��p��e��uH�憭ťz�]�3��i'�7�d�$����Vl�����A���(��N"|�3�O�);�۩If4*D�y~e	��bj�U-!Q�1���Kg�.�f����(�R��:#�!��Vv��!;�x5��6��m�݋3itV��r�-�`��\�@@̹ɷ��E��D��8�'�J�!�b�����j,ߑ#	��GͲ_>�Q��a��"�(Ä��d� �ȱ���pRi?-y̼O��c����<,�p��W�xڃ��9M��r_o�0&�3���D��#��#3|��Uu������-m��bL��]�S~!Ͼ��1��=�$��Տx#��_y���3ᜢe�}�&��]V*�4�`�Q�$M�Q~� ��i�_� $�>t������<��}�����f��sd�_p���.�P�^�
+{�m�f.�	?�{%m���3
7���)=^^a��:��^�y~�9˹�}H`�8���H��\Lc:�oY���(W����hV]xb�G�S�GTy1-o���� [�E"�}?����Q�������C8�3�-R\�$p�)������������3��fg�:���Շfe�H�����mk�`�(�C�O�rha�J���ِ��/���φ�����!V(B�P[��p۽��iN	�l�=��ఴ�Y�@�X� _dH��0�e �Z�1�A��M�~�"p�9�@z�f�����5aw�f/�07�ԐN�7#uB�[ֵ]�v��C(n����	�z� �j�fRl>ɏ�NX���G�[���dtїn�7^�4�S�k���s�X=5���?&�0�E$!ɶ��N�O�ü
6�P8�䪱Os٠ `�&E^,�mv�驻u'���F���+BѼ�[��H���T�*�w�[sQ=|&m&����e��R���,%����gu���t������_F0y�ES�1y���cN˫g�sq� ���%ׄ�`���ڱ�R�uy]��1s>���u��yO�^��ƻ�-�
�3��|3�+�>���[���W/)KbNk�G7�"V�G��r����s�����G.Ή��s��� �1��A����!��8Kҽm_�H���6^��ɺBNP��㠡�0��?C�/��&��o�޸$d3�~2��,t��0��5/��y��)I=��c��'�E:_b-��dW�VA�^���h�?���I����J O�g�-R�u���x5��lǸgT9�>�T6��m������\�a�ST�! ���a�C7�"�~m�ݭ��1���\�>�7�k��̈́'9Z��f\Y���r�������,�8���:㨭�îQ��c±M��~f+^�����${$V��0چ71l�V��PXO��4/t��#�Q���ſ���a>�ƦDoޅ�t��3T1�9��{�Qt���:��qoD�v��q�@L���pQ~+�:�k��t����4g��Q�d����N�"����B�/���rq�S�&J��`b=>���|�{%�F˴;�����%�I�P *4�����"*�L���*5W�U,~�v��bU/@rw�n�MS��Y�7�RqQn�Y��,l���@�� Z��-�Ò�6��	�����
� �W�f@�0F5M�&���[*/PrX�v�:�8�� ���gU�0H���<��,W���os��=�nskC���������Eڈ h��I~Q�@H+���t�E,"��=�nArv�;������`^������Q֝��{aK�ӰfvU��K֠u����@x<���!<�E�Ľ�%.C���d�j��R|O��7��i��z-���S$L�L�ɍ����*!B.U�ؕ�x�BU��{�3���7��~�q��H�[�=#����)�Z'��\ ��~�K>�[�);�-�&T�3���J���I���~�ښCuc�X�K��L�j�dl���J~��er�*�p��e�E����m@<��»1��'��wy�"5+r�@y�qhO�HV.Wvn��t��Э�P^�\l���ݷm�g��)A�[,�g��u]�K�KQs�*��#�X]�v]��4<���xg��H��9Ve�I��.����s��~<�S��>&"��O��c0��EL�x��m+>=�j�V��\�4���4�"�������H���G����/� c��o�Ȱ	���U����R�o�=]�������]O��L�����-Ӹ�y��T�aA9�*�TFw�s����ܔt�f���_���	�e7)���i �b������L��1������E'"�sQ�6]�dh$ /�zd����JW=#v$Lj�.�&������k�I��W�K� ��:!`r�)҇Lq�����p�=Ne��cTå۲���jH��-���@{<�i25�`�������`����\��[��w�C��K���[��h��Z]r��.ye��^�� �I�+�͖,����S$��������pFçX\�v�*�@�~�[m�����ѭ�&���$�����ڈ��8.kw����F��_$�$����{��ɐ�?��#QӰ�����g���9���7ym^��>J����$Ѹ�Sf�sy�.�sf�CRH/�?⠁�9C�s���C�1�[P��X�Ö���I�H	��Fw'��n'K���6�U��+�� �þ�9��<%�(�q��"}�s�&��C)��>� ΂QKE�������+��< |�캎U�~�-�n�X�s��B���ܸ��)���D�ȫ�8T@o�溒PW��@�}�m�7+�XJ�&�CEŦ�)�+:	�3|�	?9@��/L��>�m�ʶ�o
��:1���W�TuΏs_@wr��w���������߇�r�O�Xk��l<�R/��-<��R� 2�E�2�Im���E� .�o&X�bu�3g]��u�%:H��h���A��>:̆ɲ��9�&�E��!��i�"�����h�O�c2I��Z2�H��}�R�ݦx0�`q^X�g��x�R�lT�F�sX����z�>�K٩���Q�
X���}>�ҳ��� �10*eo�Z:�um�s�������~|Tа3�M��4�V�l߯w�+J�8:�DJ���7:/��Zļh��ڲ;Հ�m���)#ı��'������ ���@���R�Y�^�� uX	��NV��F�J+�yO�5fn#3����Ԩ��D6:#��C_*V�dyk��7��[�{1�@6�� ���_p刨�቏�^7��������D����?���f\��ff�q�n����Kg�k]�U�?�3��W�!�/C���T*�m�������`�4��F@� �#֕��o������;mok�S���*웅���h�5l��k�Ѿ��E�U5��R|��ϳT����b�Q����bT�P�"�����fӫ��H�1?����:A�(�!��a��H��ڒ�N&K�n�H�M��#�]n9��6^C�כ�,��4(��G�hɂ59�ª,�E1�4�e�=�<!S�b�l=v�.�u.�v�&��A��s�9��h\�Ώ�Z��?w���tW�f���=�zr2�ʘJ�l�d�jB�V(�(�^�E����8m.Cd�ʠȁ� l��LT)M�>�F����j8Ns���φ����~��ƙŰ�CC6>[��PF2Ǉ^��#nR�j�����AAYjޮΰ�*�p�ك-D���}F��"�@�DB$�k�_��*�Z�E`y�A4ZA1<_D�LHS��F��%�U�F�{��Cr�$M�A?7�)j�nFܞ"��|T=Z%{ az��)�H�_%&ao��b�A�����|$���=����tG�$=V�F�^��8l����k^��>�$�48G����.ͯ')͚K��F�΅?�Ȑ��o�G�?��>]5�~`xfw<��)m4�<��>�V�j�r�)�hS�t ���!MK��ƿ�S���~N���a뀙�?g�e[%���Y.�"ha}�!��^�W��N�X�G�#�x;S,JS��b���a���'�&�.nD������{�5�c����";��\�n1��ko��l#3�y�l���)e手�v-��4p?���_��L���"ɵNII$�dB^�a aV=XW��sQ�����U��5�b$��s˲�X�nc�l����PM���$�7��O� (��}�c�Z��z�^. ��c�͗�@�h��A��Oll��黔����C�S���K@�L=q�vc�f�/�Z�P�3*]�_�{�&��UOP��"tc��`�-���)�� �"���f�(uD���\�������G5p:2�Ut���f����W���`�}�a��Ļ����.	/@�*�h3���Xb'٬��X����T��=so�(��:ޭ�=e�\�(8�R���[�W����-<&x����=�Q��E6�0nK��.�m ���@������)mx[,���<��:�w�S{���L,Œ"��p���`���@�C!a�zH��)m����6��Y
�6>Y��d��4�&���ϊ�����; >|��d���^0�5�Ӓ;C��̬��vixs5���q��	��^��N��4Q�è�VX,&+lz�u�B58���秓���*5  	8B&��L�X���������ն�1���S�9��H�8��#�y]K��)h �v�1^y�>;V����x{��D��n�B��Ouq��/��|�7�`Z��>��R�p��	�H	v؏Ӑ��HI=A�r��2�(V�Ԡ�  aX&�0V*W��d�Ֆ0��"Mi���yk���	D��U��4�P(8�w��NǏ�/����aбn�~@{C��YS�_R4J > 覾Cu1b�l��{>bA%��Fl��a�����X��]{���+�n8 p��Orr��g�'���Hn�_��jߧW$��x)>V�^���ۮ?Io]�s	Rޤ-�ب"߹O����X�tƼ�3�Z$�����������=`��
��5�J������E$)�VA��d<���O5��r�3E�K�� 7��2CY���RG,�9��Q[���G��|3��ĒxKRV �;\�s�^��:��3��ϱ$Q� -)�����NG<ul�PC��q��6��ȡTK��\M����vu�Ѡ[!2ʇ��:V����9#@�EH�3_�B}�+���{ ��P��c���q 2��eY?��˵�Z&��f��x�$᷿���o��y�,�7O������|X��EO�I��$Q���u���@T$0�®B��9|vf��Գ�ԍ~��Bt�+����f�h�јJ�5ۢ�e�d2F&�o��4��T������tU76��\Za��$��,|��_ ����F�]=�u6�^���IO���Ҳ*��Y�2K�q�_�h��^�h��ƌ�9n�F�Z��E���18V ox?����8`��%�Qt�՗���4�7��0��Yg�r+Y�قn�6ǃ�SKx�#��A�f�����l��el�����b���9�L�7o��;qn��á��U-�_�T
�!�\�� i�)��s��
Ŏw��ּS��Dm@6�	̈�!���]G����?AF�+��*��2�����x�~O��g��L�>��E�%��)��F]���?��C6�s`NPF��6/8���S�ǜ^١�T��z�o�142��bmns��Z���y.�5�I7U8���/��/w���Z*$]�̼nw� 0 �i��6 E�H�My�B\v���_�```Ϯ�⶜΄��5�	�X�#���$�V�7d���ڴR�gK�?�o}E~_���~��Yi����(K�ɿ���*��\�"�!����.���˥!��(%�n���
u=�{"p�SVt��iJ*KA��~��q��TTE��p�����14$��y��@N�! ��ydi�m�ȫ7#��o�m���թ�4d�VL!���3���fhY�bc� �&g�2P�S��l�V�(c:�[��(n;K�+�w<�R��G�X<ݍR����>L��
i�Q����7�՝	3���;�����я��m�w�豫K������(>�9���X��(#���<��8��:����*��y?�5�G7,���1���Īw���°��kj�O�����3[�x��hV�.f��Zⓞ�&�5_e;�~9�O� ]����#t�l�^�
,��U����/��t�\_���0Ў/�1Z;��b/D�ANs�; 5g���Tt�qQ��$�2���l�#[��0H�Dz}���P�|�V,�$J3�=��'EŒ����]�p��И�^w��`@Kc!1۳�P�Θ+��	O�el6n��]��_dP��&��K5i�A��ˢ:��5�kkK�m&�3�	Jv�5{�� i��]
��Э��&��q(�'�n��MdR�N��緰=��Ź@G���G�wE��`��T5=�X� �<� �=0l�U�(��|M�D,g�/q�5I�qغ����p�0S��\�e��_{�1lp�l}�; ³5.�����gX�6ȹބ�g�sO��|�lϻ�S���^Ok,���>2�1Z%���YT���\��g��"*E����^ꊼ�͙0��S{�󏥵�E��K|�'��)�{>��1��9/��$M@=.?�u����7rRz�3^�씳���˭[��F(���M��V�A[�re��:����6��7k���g�c�.4�Yľ�Jv����J��⿅�c#������B�X�[�C��Q��'=a�<PO���J��;2U�X�OU�سݿ6Bخ�In����>�8{׻g-՟�95 ���FקH��('.��O�&��$y�o
�w�L��ϸ��"H�J�N��)�_-�\0�'��2rO��b�nuv&t�D����4r!~bj�7�U��>ƤI�X�7E ����]���إ�Jn��݉�\���ǋ��4d>�#��\ť��h��/��3k'��	Ma!<��k�l9�K�%�M�/2�i䴾�FǺI�͊��A�W%3����ݵe�$��N�`�aa����7���0�������:���4�~�Ȩ9 y2��:���Q��D��l�lA-l�N�G��J�D��SYw��klBL�np�,a M�*����_!˳qI�0h����}�C1|�����?SY�dq��T�k�c�^c�Z�P�v<��l��U���R���A�%�������։4�r:�+��'�n�8ϓf���ۻ\�-O�����K�Wq�s��$��d�D�+x.��:�˟H�nQ�'�Ɵ� ]�/�|��9w�ӕ��h��V���/|���7N^�6ILBO�e����ۃL*C� ��lЭ���E�+�Y�&�k쵺c�$n2�!}�֡��b�������%i'���6a��Ы�8��ݛO-b��\��u?��l�M���4
Lq��,4�Ճ,E�oF~t����S����(S�5$"�,�C��ڡ�҆�<;�u|s4����u׳�r�읭\�q�E�x	`�ы3%����!2��S�)�.�����H�1��R0:� �ra�����&4��	9@���QT�K������!xPzN瞸���,<��w\�G�t�&?:eqQ/��iEg6B��CLϕ|!����Yp�3��?jc��F+m�]"F{��wCp[��^=��;���N��nN��Q�+������U�E	>/�5�Ak<ڳ���k�M��@����Syd�#\��7�,w�pS�D�po���3���S�����F���{�d�#��d�s��w�?���.e@�m\׬Q�M:�)�&�z�jg�]��f�O�B�S��C��z��̨�kNSZ�K�a�CQ��e���A ��D�`�X��4?R0�4�
��[��VM·�?���LS���R3�Tٔ�f�0=<͍S�-��E�/�F�wvo�b_�"��v, ����c�ü�]=,sUj�M����h3�YO��ܓ�=P�H[�7;�{h�Kc��^{��SH���v �ܗ�Ϟ�}Y�>,�p��D�A-�٩iI�g^�S=�������R8k��_I7;}�JL�����k�ո�
-6X�0[��>���a_}mI!0�;2٪q*�"Ǧ���}t��D0�boI'W1�W��=�?9�פ�ɶN�G&:v.|Ob�Sc�(�R��ʪ�n S"%h
2E���	!ˋ��AE�d;�P�C��gg�1}�f��^�&�F��-�D������I�	q��lY�%��&�,��qx~M���綰j��AW#�xF�5 \��w�h��-Q��U�e�-�3��Y4����΂�G9���
����tV�~�;�u�8xL��`z8��l�%}Pc�(l��Ŭ���uvA�lx�啗�,��QIC�?��� H��P}8��	Z��\�e/> ��7�tb~�ˈN_>�}�q�3نvT���f$��S;õ������"3N5��e���8 �?",�y���Km m���(C�����_,��g��
��O�ܳ>x,���ﰢ��0�	��� �xo,+�7��[w�z8�(���g���ҕ��$����([u�Ů�e`F��W�H�%�P�e`,�B�@�-���L��s:��Os8{���o{�<�ͧ�g���R����6��AG!��F'H`��n�uj�$�EO�	Vb��9K0�۲�(<�.2��c�"���� �~!���E�Q�� Z�>�oh�[b@�������gA�H)ڨ�& ��x��._Й�C�1hi7A�xV����G�W�����7j���m{s����Z�:��>y�w��/���o�:��G���^9�7`��<�(�љh�4���N�r��1!�uJ�O�b��\��&b��#Hλ.���Gtʯ>�0&�1'�
�
��,��ή�H@�ޢ�t�|������Z%���t�OCM��ҏ��:=W�햖R)��kk�0�@a������l�!�h�N?��;�zB��ۚQO,Y7�H�%B���f`63�m'�dp�6�-�O���UG1�} G�&�W��#�4����+&e�#���K�&R|ƺ�t�c��sk`��Z6���WĊ*�5ʦ���]@�wxm��,��h.>���.FŚđ�1I/�6����J�Ng@���_�4�����#V��1��p�37���ˠV��ѣgiJ�)f�\�ʶ4�Ch�U�Q������r�r0p-�9{o��(��'������Y�XE�Yq�&���ڲ^a�[פA�;���w,�cY:�ɋ���@��T�1n�`}�ӞVy�P��7o���~����s3ǌunA T���,׸�u������N�%ؚ�{\3�Ì�h~m��C��Gh�)!l��5 U����9�w�	�~�sR��b��M%�6�J���-�C����FS_�-DqO\K�3�:)þ�sQ(����z�����k��_#1�i8��dh�qdy~*�9C6Y����)iq�M�������Ü�)�&���!��<}R3��Jkv%-����]�YE֜n?�e��V���.��� �t�[ �cy;$I+��)�H��T|�*�y��ţ���0E'��i��m����2fV�ryL�����
�s] x������\�
�� 6X8TT`�����e�`A��(Im��3׾����5�(Q|��T6��"Z�>T�HT�x��F����#��0�A�_��_8�ㅨ��TV�u|3_�b��0=0�e��@��X���鶂p��@kWmd�tP��/}�|�N�]�?Hܠ���Xn��R�L�;E�)�tn<�#����pc�aNL�������I?/O�x{*L I쨾��s��<܀�)�~EA�j�t�����Hu�:u̇��a�qa�
����s(4�1L���4�,��5y*B�FЗ#̓����B�`� ��Li�.j�����\U���;��l���N�]�	Е/�nl���-0f�m���>�ӊLsU�;.7�-�I=��.GE���6�MT���!���������*31�
m�7_v<W��h�p��2� ym����p��=�'��M}�<��ʥ}ϏA�%2Vm-�
�j���ȓ����H���˙�ꂉ��%z^� ��ob 	��2z�l̓5B�5b���3y ��Մo�����K�}����Է&�4_|�J��u�`�S���yf����Z�R�!�<?_�jo�	�V4���B��&��Լ���MF��S f��O��0�z�����w��N$;5�?0�L{�5��h�R�\/������X�K]C�͹���|��櫹��W���İ/#����%���ׁ�z\`�*����O�3���� �8K!�?C\���!���'�;��C|FH���kj�G~]f��n2��J��ސ��AY�I62�@�6o)�V;`��>��:�=���=�#�5�0�Vt��4Mh�h�vQ�IQ������nm��ܘcMoh觖ېK���~��Wy
���`���bV
%�����g�f�3p�,��:�iN�?k}e�sЮn識g�r�[5����̲�r��bEm8����O�n�w���nA�V�$�`������d3h�u"'�ioB��5��:��RT�u�Nˏ�¥ƍZ�D�k�����bEN�4 �r�k?�����p7q�ÜVs_�`����c�K�&�����>�b%�P"��:�L��zt T�����ǣf�� N
�BU��U���Q!j�.^�ո����: ����rؤ��[�A�����|��d�s#�f#m9:_?�u9A��l`=�H
����>J�����ϐbI����2trHD��n�E��M銧FCZ��)�%j� �7Vܜ��$G{��U0y߱����e���'h�?M���	�H��
���� ݼƕG]ն��}����m��t��M"�{�W�e�=��(�N`��5r3z�K�N&��7��]�B�8+�3���Å��V�*n|�� �G:.�� T�8�{�����*����I���PL����)+�h^�XVa�l�@@лQ,m?�%��L�[�'$���ܲ��Ur��&��}l���L�Ȳ��\?��dT�IS����>߿-��9�7���\���nF�_�H�&���v�W�ez}U��Y2�vҁqA6�w���3%�٫�^�S+���>�q��qZ�r���~H͗�ڡg���A(����`x�s�g��(ؔ�g��d�8�p���M��U�7�ɟ�������X�.�i��ծ���|5sQ�U%p�o-c��21����p�8�`
|�'P���;t��Q�rf�Fa����?>� }*��I��,K��znN���9M��0����̙p��|5�NIQ�cP�崋
0e?�IY��U�A^9��֐e�3<={��F�s����oŹ� I�)�Sɝ����rx�C{z�A/A�$�5��V�q9���X���*���d��� �Ւ����TN���Pw���D&i�P�R�$�����}H���V���/��a~�X@­�τ��̲=κ���Q�)\�:�Hwlό�b�����9�\7��gT��B��hz�w2^9r:%�>#5�!/�%�al�Z��/�-�p���.������,��h�>!abM��q���hBZ��T�{��/R�`�N�a���yDBή��N��4%�EF�t9�I��9|��Ya��@*S�o�>QvO�C�� /�_{JL���X��7m{�X�,{�ȶ����?n�Ē�� ��XD�P��!P�*��C���n6��y
y�-�dX���0\Ky�~g�j>��xP�B�2l�r��v�E���kD�c��67E�-�ktТ��B���Xڭ���������L�Mo��xb��+��n��'��Y�����42ߤ�!�"�sO����f��yq��YQ�$[�Q��~&�v4���i�f�w�z�\�]#�ˢ6ۯ]}?����e �h1.h'�4�D(�f�]�"�<�`�����z5�SH,��$�]���Y7�-&�~����UK?(������(vP,� 	^4g�*���j?J�t$��"6T���^���chɶ>s��~!���iQc\�)v1Q�5�xP2�~y�eR���Da�͹_���*�:΄��w3�<�m�RWfLb��C��#��qX��I��9ڋ��V����
>���I˞XE��O�͖u-RD6�c&l�el=y�Y��ۧJfvs���&�O�T/�����2�xs� ��Y*��d�(�s�D�J����gN8/��H������h�Bq�+ߝ8�D�X�̢&�S�Mwg�%���տ{0��Ψ.Q�N̹Q��O�$\�c�?�@:����刟�8�Q��8v�O�#2G��`,�h��Ҿ��s�CX+��7��dv�79cV�5u���Q)6��'�v�lm��n�:%�v�x��5!x��6���6��A�(M���u[y����d�8�_k�N�>���o���%��T
Z�UP��'�-�ZU�4.	|
v��0Ϙٺ�R�Vp�t;p����m)}�$�x�Y(��h2�֔�`�*I�$����kd��G]��E��MK��Tl�M�/�Gd	DC�Ca$����ŲP5�#3k&���_r���;ax�3��F)t�y
7xN���KTZ�APX�/���vОd!֕��̗����Ր1��+	k��ͦ(<��o��*Κ�=�W%���%�Z��*��^��.�b?�1�ؒQp��E�N�b���c �9#*�hjwl��G�
m�QO�����
1�|�.���l���7Ԟ}uP��}�r1f�ٷY���r_�%3�;�Ք���s ����]§g�H�$��d��U�����v�����YD2�QIL!�OΏ�8�+����燱T^�`@�8��������:�c��o�!g��Ϊ���r@j��f�%X׌u�?S�T��z�z q�ʞ�9y�2�
NvM�F���]��7��>�����މD�M:X���*U��~x�;�kR��[��E��* 7|7�x���7�GU��KIRg��-�R����ؠk�^ymCb���u[���,kAD4O�O5��m�s(7�;"'�e�	�b^t^�^V܎�(��St��D�J��Я- (C�������Ȕ����oj�i�J����\���]KH7��[��N;�`Lm����\�,��IPʦ<��a�|&;���k�Qi�ӣ� �2����V�._��:��5�T\Je�eХ�m̗yjx��4��T%侭H�q�6�7���՞nqH��<Զ�I)-��W��wQҎVq�..0.�p^��н^�~�<�틴��G�2¾6����5	�"�b�܎��e��ƹ�&=����ȎO6{�r 4xi�X?������f9$ܷ��˳��j���\�W�\ }
ݿ5l�|��
<��Hs���u�+4� E������A��M
�����$F�tۊ]�-���˦���$p�榞L��S�:����W��h@��,5���TA�Sm�d ��w<�C�FډX�+�U�G����U���ߙ��5G�Ƒ`�eZ�s�Y>���:�	��p�^��J��,E�ݪp�Ⱥ)� �N�`Q�t��3�0�F�rF�*:����~B'��)���^���4���r!����5ƴ��	Pd4�BR�wB�e�)1;S4�ߴ���q��~}����{���r�v�wďع_�T�y�Ő���E���~��%5`����}B�{f�-2�����$�\4D����NJ�f��dδ_�-ս/�B�^`��Tz�`�<Wh7|g����\������"�j�d!7��2Gr�!t_K�.�����^o������q�u��\\Wn$=1�+3I�Ř���r̨�d-��Y^p������]���$ٸ��#Sab�C���
�$���ݽ3 ���dc%Q�
|��A�~�
<��$jA,%�?m�m��B��=X��L8�#�y���b�ei.�[Xm�<-JR.s���>�_mr����Ai$p�G�zJ��ܡ'Q��?MS��iu�k#�d*<�]����� �����oa�}rڧ1(��I��mڏ�w�0�Z~@\�D�-�>8uڿ���$��Y���LTC�[�)S��@ʉ��5�����	t���u�d(p�����i��n���^lS�R.dR�N��ܼ�G�'P���Jk+��Mt�냌mPdM^Rz��P�T�b!�qR��7r0Al8�JlL<nǧ�(�
�A�hU����C��O��A�4� |T?���'߇%�.4��5ݲ7�R�!�e(ji4��S��m�D�-�~>�2\�,���P^���讙����R�MŽ����M~��˶��B�.���%�}�����֍j������eO��0�k��̌�[��n���i(/���~��t�[͸��)��Gڡ�����!����}����C�H>Zޖx-�$]]���8�
KXԎu�3�E�@��`͟�
�N�F^ɲ��Dt�L3r:aHI�;��� ^��{^MR��M���:&߾��Ǿ�T
�9��c��G�NL��-����%f��)�k��(Gبr�8���5J�� ;@|�ͬ}7���!�|j8�M�����ʷR���x�%}b��h_C^�[��N�܀����\�����sU^�qK�2Xsj�~���j�y�� ��+.y��NY��l:�)�gP���m=���ԙ���8�]��?��3�r�)�t�/��E	<�ƺ|r�`����'O��/{)�'�gh��~ȷ ��L�:ܙF�*��@Lr��t����h�D���zX����� �H�o��N��UR\]*�~�*���ѪWw����B2w���W���W�p=@���{�}�,�����Z�K�J�`K�� �!���XG���?7{�6�c�kgD䯠��A�fy��H�dC��v�t�?��$�lhC��pCfZ��Ae�Jҝ.}8��Fi��	���f\�\�nR�B�\����Q�3��X��D(���v8�����pq�Yt7��ܐL�p,ʇ폄���5��&޶~�Y����g#)K,%����9�;,B��|d�'�!u.W�;T}�p����bS9�X�{�P�K�P�� F�ɽ�����5JQ��`�7?QP�]�F�Ϯ���NDz�Cm[�[�f+*����O��6A�-�ϓU�B�0f����	�b�`e]������'����VOF�\8�������7�m�o^H��u�L�#j֏P�#��E��og��z�vl�W�j�0(��kl���lǴ�,�B�R�ށȈu����j����P�q���Tlݷ�kKw=��BD��@Hwj�8�8�}-������ⰻu���Ƈ�^��Yʡ��*��w��*dd���k��o�C�� (+������A�UQq���{�7�|�d��S�z��S���x��p�q�<���q������N��r��9��N�&�V�6]��1
9z�M��¸dX�������MI߮�"G-�|�)qV���vH�>�fees��ig7�qW:�|��Rq�mQ���s��&�\ZV����Ѹ ��P��r�+��F͝V/.��/�F���ˎv�@�u�"�u�x�rM��ҽ��
�S�`�7~2�̤wK���Md�y�azK�Z��Ƚf�����~����d�΂��8	Ga����ܴ���t�VVG�n3 ���m�s^�����L��м��O�\yC�/����M�<Wr���D� �k�[
׈����<-���o���.1�����<"2W3�\2>�1��m�4=�ѹnkʾ��T��bZ�� �-_���������r��aϚ�1N�4�bC�f�җ���ek��'T:U�X�-����Zq�#g�a�ג	����C
�t^���Y|�[Kl�z�V��pԄ��l�__Ӌ��e�"[�մ��Lv�Bs�Ũs˱f,QB�l��tO�ZJ!�	�{�s����g�T��Y��^˧�L���7L�`{I>��2�ڢ.0�rB�oZ��R���.r����̢��R<��y���^���s�Q�S^�����c��?0�'y�Avq��|;�q��������:HQп���&��J*���N�]���k}&��G���d�n]�
��RوP�������N�p!)����W�W��ʫ ���<[:2���*��uw�&�b{y��rB_�^;D0���E9Zw:}�L��"ڱ-��2b�&"6���O�j~N#��25/��Շɟߐ��X��=r/�~�q75y��)P���@�n�����b�w`$�lϹ{�&���2�`���+��Ɲ�?R*���p,aI��5�7�c Dn�<M�1�"��l6�WWO�˱�ҥ2wa.�<�q<����^D���LM��t�w���1�D�F�TO|uCw�~�tj�/����a�]��E'��F�Z�`��3��E��77��������Ȟތ_��"u�M�V�?h�#��Y��w�R�Ŭ
lͦ�,r��N� 1J�"\,�J_��
��s�+^2�?i�L�8�K�� �� �_F���[-�����3�C�/\m;�K@ՙ.O�����~��fi���dI��u��I�����/��ٮ%�Z&eI-���0�d������h�u�������^z!�l�'x;�e�3�|��8�^	��~�4l]��������l�� ������<�-��gl���f��$��s�u�x������QRZ�s9�Ќ����O�Qj	�͒�gPs���a-w*��Z�����F ��{~B�L�ɍ6a�;]�*�i�'��~U*�Im�����C�mT�\�r
,���7>���'��0W�]�գ����hʱ��l��>���]�.&�g{�P��:�OTe�& E����Q��|R�9䥣� ��ޯ��x7&0qUf����� �*����^�a�$9έKIг8��I�.�Hd�.�S���}7)*��6=RSn��D��5�}�E�.u��Im}9v��H�Pb9�����\64�"mX˖�x	?)�Hk�ES��ۊ�]�H앑�?�� �9#4�}���	����Hއ���?��S����P[�mk��*n���S	��$G�V�Ŕ/M?^ߑ�Gd��)\��l�=������GU�+J�|%�=ۤ��G�8!DE<��pQ�k��@Q�)�����p����i�kN(p",$i�R��5��A�Q�O�H#˻�<-�V<;�U���)�d�Ȋ��刑�i$n�8O�ɤl�V�Es��Q�C����^����mn^*?��TK<�� �dpz������L(EO�6� �߽��.�?�n�X}��p���{�_κ�O6	���ϲ]ڃ�*;�må��ゟ�����5���n���6ң���ã�b�r�V3� �-VMÜA�ﯧ�����l{+eP����=0�Ajta���˅{C�u�C�Q;"\�[?��_}K�z�D�t�������`f�0M���NhW����$z�j�_"5fI�w�PW�_�Qs��$�����LLWT*�3SMv�۷*���/��Jo�]��\X�>\�~�Q��v7%�����Z �<Ni���[��V(��,���A?�J�"Sf�*�P�e��Î�́Ī����<ͩB�0����<���5�3A�~�T�YFE[2�dUْj���S�%w*�h��ӝa�[:U�'Rвi诩��p>P}"J�%j���O,g�ܩ	�b�\W�k��)OO9��}$6����)���
Ƅ��2�In�+k��	�k|��k6����Z�Uc���1nn�|�\	I;�ѧ+��s �f��������J�z��q'�Ib�R��ܲy�P�m:W
�û���nю�k�M��Ei�:}���+'����]rC���x�)NtW�t�5��$�����2�j�Bv��u,Ą���'��0�û����au�U��S�Z��>�c<�V>�Ud�^�(;X�#}̦�;��?˅�`{A>����.�7�^��l��U.���	tb�$A8��'sf��J����b�N:�bEn�y��b���?�}��;dM������;��T�~�.���_�m��1f(vl�x2\��P��>��l�t1]4ok��(B�P5����Qޑ�E�}CX^e�'(�/��vܵ���&V�aW�&a�h��es�T^�9�L�T�������;��`��؁�R�(�Q�R�P63�� �W���ڠ�7O�����i��z!�?��S���F��Q���A5TI�y+7o�Y��:^ց�<��
JF�󜔳	��mϚ�Z	�)L����C�yg�ӧ+|���7.(�Kj��a�I�Vz���w+��ٱV4���1Lƙ��%4��0c5�Ԝ�m(��R[;?n*��O�kL�d�S�	���_�M�%щ`3�N(��C��h��T�Y�mo�x��{-�/}wt����ǻQ�z���Y�k?8U�K�
��bM�:X���l'�j�L&�/BJ�"�E=���ك���\l���!�����|@&hJ�2��Sਇ~�G��C���S���%���������6Y�K�i����O���u���W�K.�m[�3��|�&c��ŕ�7�Ϗ�JM�X����P�m��ۈ>*�����܌�1$��^�~\�D�TG)n��wL�z6��D�l��-���y��ۗ�/���;��nN�p�BL(����X�'��i
Ŕs�B��Er�mIUD�@�a����÷xh==���E �
���7_"�|���q��{���C hܹR�QZ�M��n�gG®s�'gվ����9�}���j)����l�*�]gSr�#{�b�U����� P��������Qlƞ�
-�l���<�	���	>>��~���g�,���m`�B\�=�y��#�Ef�;%�>���.�`�o�+_w�����dP��_H-$�?��Q?���joć�9���,L�D�\;�X������Տ,����[4�U�$���7_1�J� �QY��DUXX@���W�mY�Dg�.�~o+tb{������#�vR������:�x��29+�[Ѭ���a�UƪJl�Zʛ�2�[O�I�i�:��c�Mű���x�d�1�p,�-�[2#�b)|t���Z�nm'` T�ڄ��i����Sժ��v�����`�$��|ǣz[?r�8�XL�ڐt���ڳ����!Js��+�h��tf�F��?� �12F|?�V�9)Z�`)�����t�so�\�0�m��lI-^Z�f�X�`#�	l�R��A�����Px�4 isd*�4eO�*�l���Ⱥ[n&�����BРn+�����j�)c_�L�`DF�`�w�.�?hxĶ`���v�,;��!���|}��B{��hH�RH՞�~o�F����*�D[�A��i�e��i�"���ҲF/��mLx�MkG�ɳ�:~��>P!�O3���]S`_6=�G�=?딀J��C)Y����c7��'͍����GKX=����m��Y���ޭ��D�-~F���I�C��;Vp@cZ.������K.��%s�:)������CZ��DV��e����0��*"��2�Ԭ��~s�*d����\1��J25L�'���!'����/�ɪ'�xb���{|B�������O�;��\����m��rᷴ���y�᳨C�������?昁�y��o���7w�Mi*��z�w՝�&���p�H\��<���&����R
߲�E=W�܃V衱~�h��Ĭ��	bS�<\a�m��Q���̃
t%Q�:R�uOH�I�����U���z�sa�j
 �����9��נ�d ��l��"23��ڿ:"G�a��<���L�f+!�(��L�\,\����]YG�a��׾B"}�[���p˒V-�. ��^�����A�{�b ��S4}����P�^�0` 8a���.t�|��C4E�"}�����b�#�#��K�ba������m�ZLYD����%�<�N���r��Nd�Gz�L��^���z{@����ؘ֒N��'/b���K=�j�?_(2�$-}�.�������^���i�T%9��B��f���Ea3ÖyEx��Uj��	R�զ�n�Dr����� ���瀞�OU�b��OA|ğZ��a(X��'�"�!y��(��Vj>>	V ?������<�G���ͷ�اK ���<B�߆sn�*<�����Q��z1l>^�����Jk��׺H/MS�#�����$�#���Gg�b�zD�ݎ�m9�$$K��ے�UP�dy(�٠�������Ĭ�|/d�.a�T=|?�S��_袼5%d���<e�P)���SUk�]B�Ѧ\�W��^�P���@�bQ��bf���,V��ASB��c�M,�"Sn�t��im�+�3-�Hqwش]����+f.�{�7�B<�S�i'@`au����yP�K k�p��v�k�r��2��S�O�Qd�e|�&�ӥD�������v���Qk�i�P��HqC�\ƺS���x����?��f;Q���m��m̲k@�*9�o�Ǘ����ז��I9��w�H_���YT1ȇ�vz�\�pN�V���Ǭȣ�Jw��o4T�N�ւn�.L��[^�9c�ד�1k�ly!��5pʪ}+���܋q�7+�8&�����<N�K&�=�&�9T��^��Эc)�©=9�')�$Y�Ύ�>�5���a+D�]3O�"����+�Lhu����t�Ꝺd��E�8��{��K��1@�b�g2��]��+�AdP]�r����hi ɦ݉�m���Zևو��	�.�1���x5�@�%��|ЂI�_!��ч��9,��c�F(�Ø���FQ�T
I�22K�֦�a�G:�b��yY��F��hh�7���
ph%�03�ng�+�����(>�[�g����rkG�)�1a��W{����jr��?�-���)�?�����N����ba��ش�)_ؕc�`�\����|/�Uh�2�qr ��;�Q��\�<~Y�����^RC,ϊ��Pn0�����I=׭����*n�;�����a��S��j3�☬���
j�Du35ڕ��ś��	��N���U���V ������>�8K��4�/���6�������a	S�T���n-�� Ny�CB�X�Gݧ�P����D�e.1�]�3\;�>�\�E���f�0�b7�/y<ϛ.�ΣB�@�(�L�� 7�
�Kz/�#U�R���*���,A�Ҩ�o�<?��d���O��ō+|Г�y$���]q_�r�>���գnTD������M�V����U�N�>����0�	T�y�d���?����yH�k���p�2�Y�=�(4��}�A��yO|���(X7}����ʊ���J2��F�B��[���W���)F�&���&9˙u����9ߴ�����1�7u7�8r� ��0�N�Y�n��*Q�I��7�L~3�1��,�	Xy����Y�#Aw<E��`���V��x��eW�<����U�:���b���Ɠ�r-�<� �.W�E&�T�I��Ŗe|�Vy}J��F�E�?���|}�&�.�(��� P���f �Y��4B�����N
�;��e�]"��uPתC��	-�x����)<<�����C���m����4�|;:�>�n$�)1"�6d�g	���bnߒg"�u3�5�k(=��f~�,�p�_y�"�:�Y����1��
�k�	l>�G{�p�}�`״�,jH�n�`8�#�q
���h��j-�?�Fd�^��0$�x�KG��5�'�t#&/�≗�[�L��x���I�� ]��>��>��X��E���k+<�:��aV�q��c�r?KvcQ�h�J�<`���M�6�:^�������&EQ�O�D\`���^��P6R7�ё�O��%��j� ��+���FTkV͖��'��5;�w��y�V�!DYo��� *��OCj**��܏���A<Ե��,��׻�}oF��
[��%!0}E6�u�2�B���]
1��u�p���N\��u<DF¿��q��*���D]�q���ԉ����m�i
Ol�2�P
v�(��m y���{Sh#���H�l�.�%�#b���]��Ull�=��a�FzJ��Lʔw�Bz��@4S�V�jU��SŮ�wq�K=�_Ckrmn�
&zh��uCe�*�����]R5���pG�)��I��������^�hg���h]��"�=Q�M�l�u�#���[��ZgC#	�㍧
#��S��]���xj�	�EC|d�]lB.X����������a[��?��ҧ�&(?���������/N^[��,�j�W�1�������e?Ga��7�$ypO��)� �F�����<_�x�B�捚eU�}�sH��d�+?��xM:�]��Hj�I
J�`�(]\�Ǔ��ٻ?��z�����3�J}H��?<l��?����.�wywY���� u�J�� |�뿒���O�z�[|� ��3:
�2� ���6 IS�ٯ��W���E��_���!���� ���(u*�����sJ}r��1eAf�~�dr����eJ�)��j�낫��q�s�OYũ���	\������Xӵ����|A3C*߽W�0t�m�ؼ���ԙ\co��.p�n>�)��|�^@;/�?�	xJa�A$��&�w��a��O�t�@�{�e�d���	� M���]f7����{#52<�SE�3������E�6`���bg֮�導3+)�%~���_��1�3�`E�v*�vC��Mv0&��uMY!�/q
���3�=t�7=��Yv|L����uH9�w%��K蝹�Ya����؃��낖z$�0����U�=}Ff�f֗����ז�oX���6�˸ڬ��OyN5�!�������5�;��L%��{����+���yE��èx�"���U��E?�������T#w>cc��>y;��&�a��N��`��}��d T�}2����u<�-߁4\@b��m�(��̬��?�� x���Jxg(^��#�,ң�H{�����ڀ�� �:�Jd����$Qi�4�4�;�~���o=��RVX��8�O9�l��,7�s컎WOȹ	<,������r�����wYS�a�÷9�hGIl.��ʣ<fd��K�=��	��b��꽠�����]!��Ӓr2L!�ʽ�z�]�죯Oh59��(���o�/��/q>��񧾄mN����j7N+ظ���Ą�������)�����]��*�R�Ƹ]��Q��Ϊ�L,㙓^������F;�U��BP��-/r�ZY��}��vm^�]���A�gF^��g9ޣ�=  !�0T�*�N�`a.���?Ee�r��}K��R�W�OH��� ��Ʃ\ǚ �J�De�ݷs��B�Y�TH���6�>B�dC�޷�9BDB�f�U�'�LW�@� ��m��L��<��^�i�����Ȇ���1�^W��&�$Ŗ�����xc��3���uJ¾W2�yq�vZ�P�����mW肰B��ö�k�G	����a�o��D�V�T�*�W/<Z�� |��gϸ�l 5|!�0�ŵ%�5x7�o!�YFR����N��x�a�6b��3�?��^LOPN�L�lP��*}S�Xs��tk�#����nU��M�� S����Ⱦ��_ǌi�^��v-B� �W	d���P�z|�B��)'Qr�|Mׁ�:����gk<=]{�'`�ƑC,�F(�o�&~ѓ�S��(�y�ݸ8k5�M
�I1���a�����Ǵw<�������t�ř�c��"����%7�f�+��9���<�n� �|ɣD� ��i��#đ0�Hv+�釓����]NZ��Y���_3 _��C֣��m7&�<�b�T�U�3t{	2�e%�l�\O ���
�è�6��'��_��b�����1�����co!N�z��0"aល �7�(��p�y� �l���~�̓
%&]�n���S#�X�'	�	+�Q�`	��H���P-�
ؑ��8��#��_�$���7x���Ct���'.�-K�c�pOݘ�,��.�F%d/}����:,w!	�vվ:�����@�%�Mh����,1W�&i"/���lz�w^G��S��}�)�C�G�Rn�XJ�<�O�ҹiN;�DÞ^�:��qL�m�v���@�SO��#?�����Y�������	@�8��J�QE@O�G+�V���l�eA!)d�Q�xoI��$�0Ut�a")����ۦ�)� �w����P�)F�Y�#� �{���I��P��������~]��Ka�����ӏ1�.�OLѵA�b�R˺���d�����)��D�>�X/}�4�.���(*��R�x޴n�I`�2���ɽ3��4&��k��x��Z�'��]ks.��+x H�1�oL���U���� ��C4w%z*s8���2$�U=u{v#-�9��:Ѩ:פ	�MhU:��G�gS���-���am�WF�N���S��O�"R{@[F{�q�|���)��P�oVa��;Sm�a��y+�����)6�s3���r|3vܦ�/B4����5��5���g(w�ʟH,�8㢦j�6��7%��_��:e1V�-.<Y�'3Cek���a�T��r��z��'�ܾ��Ѥ��P�1qR�I:e�ו��y�%lANe�<�[������`8׍6�~�va���g�u��PsO�f�W�"]�+���n�_t�ɈF�n�iCw� �D��>l��� z��)v���0g�!�z�M7FQhv	K	z>�2��n�.8�e���WI��<��ÊA����e�6«9�����������O�!��Ŷ�m���w�y�i�4��YCSF��~�x�U>�!L��]g�� �5�e����RV�Ԃ��6�U�B?l$�/���P �W� ����+�s�>lM�G���K�9G��T�Ԟ�}����x4��߾����U�<���ި��&�Á�h�i`�~fǰV7���OO¸�6z~���*q-��������4Ԃ�uoQ��u�d��h�O�$_u�\]��� ��<��&��'�3�W��f���<l�fv���	]�X�&֩&����+F� N�T�.�/����f�1�C�Őg�wkT�]�s$�F �t�}���C�$�įc>��y�y���>���ldq������?+`���*3�]�6�׾)�r_~�I{�a���,z�3�Bo͏���qM#иq=�r�����#�/�O8�<���`}��qaɮ�=f=���J�����S�;Q�6~��Sŋ���Iؚ�Z)zE��%���	C�?6A����k��ye��7�GNG��L��C�y��^'���� ��0��'�����2�h|k��(ՇNn��ҭG��u�,<L����:iT�R�np�r�!ѹ�GQ��5Ȱ���7D\^�i�Rpx�i5������Î����B�@~���78+��{\����m/��k+�|Qv��70vb)�Qh3�:��2��"b���hXڀS�:��~nE*ūtI���Ǽ�VV�ڪ��`���č�נ?0���ݻ��F7���N�!<�'���ZOcI�?�{@ߞ#�ࠑU���~gx��<�+�qX�
�r0 �3���Ə���L<��6)��ny�{��71��Nc�������!��Q��{���G��Ӏ.;e8p��}�D���% knoo�e�1�u�󖠞�6
Ac���dfS�"�f��e`z	�з��/cT���ښe�2���%����$���K����ɡ`~�	]s:���$.i�4�ѝkQj�4�qb�H��A�����*u�db�x��� ��P��kc���y�9��I}���s:+�3��_���8������/o�oB5Gn���z�x������zJ�!��[��S>�՘���t�6M@�,�*�e�U�~JcfE����9K\��Ӗ�+k�:�ɕ�^�,��!i�������J%�5Tv�ؔGB(
VW��yl`_����?���H_�v��_���d��aX����:m=�Ǌ����>竏����a�é�v�NI����r�B<Q�ʺ����}����Fo�=�T��\�Os�p��;1���9�C`q�e���XV:؜�FA��m��eO��}?4��N�jIU�F�i�M���̣f��N�OBX�Ol���7p� UI���8'sdGΟ�7v@�ص���ė��.��^؎"����J�k�) n%ѿ��!�dn�MbW����"�zF4*=�q9�cĭ	�>�p��nD�u
[��kj�@�:�,{g��;�<wWb61p�UW/_��H��e����H-=�P�d�|HZ����n�H#�J�_ċ�?�b3;�w���R���@A�d��:W�fT��j�A-��@ģ|h��7��)5B�J��|�4~�07K08�ś�Lv���Q�Чrڶ:���ƺt�(��ȑ�z�u>���/���oZ�|d��d�@]t>rnH<�VU�ճYgкbN��3F�j�@�G�)dK�x���̍��mo�bD��,��c�.�MǛ=�\QZ1��L	=���XCLZ��QeƢʠ��b
���p�p��xUt�c�9�3J0��~�:�Ov��	Oqf@d�����aϹ��X9a���So}d��8u��,M(����9���`�������d�w��*��a5�u��8x�d��.
��᳽`��K�-�j
}/dnYoJ�0�gL�_q�ZÏ����>��@�ii�R��3�xaLH��������/i�Ҭ?爳��l��'�<���$�g�m4����d�:?��������"�	a^Z?&Y��=����.�2'�K� ��B���!��3L0��bBS���h���C<�]��n�q����Y����P�X�w���z��JS��4�s��� K�ݕ�0ʰ4UeWE��}�z:�:<[?㦻 ��#�Tg]�9+Q�/+�/�q���T���������E���p��y9@�֖M��Z�4y7�m�.I�k��Sp�ȿ��9�1���
Y�p֑��〭�3sAz,�����9�x^����pe�J�P�q�� ; /�g8�r�-�q��@,�6����Q2₍�X��.��Mb���3��U�?81z	�;u�*%���Ay��|�ۈ̭��\dQ�m@�$�!����֓�޵R�#�]�\��4=IG<�2B�x9�	����a<��+��a�)P�J"rp�{����.&�5�� 8���Y�O�K=�F#kX�V�����1�M�KB���1�Q�Z�_!�2G�7Q�(8H4�5y��'�K���"�� �;���y�� �X����kJ��"g�%t�y��=~�쿄sD	5��[�.���YZɫ\D�Ǟ#Kc�z�8*�z�.�me�^	&�����)._��_�hpS��B�j��k�'����,�7^C��"#�1�5�~$���bd�`�C(�����d�X<)BG3�kO��8Q�]�![5���xr[!�ԧ��֮�<��_L��]ض݌u5W�x���c'����>A]����g�vj�n_����I�����,s��>k+�۟/n�����:���D�|W��*�%�l����m�(�i�[N��$�ۺ�b���vm$�'*'�a���!O�^�ED6�T�L��>�.	f�Զ����xK�Lh.��,���eZ.��y�: �|��P^،��g�s���e;�O�w�[���x��DV�Ś�P��ԆVe���"��[��i�՞Kz��_��Т�-'�������.���܋R_��4���� L��UE����d�T��\�[�4C,�� = ���]=2�~0����Q>���H��L��3�leLW��E8f��!���4���*?�ln�H��n��p���dY�D�����wq�����(�m��tv�y�u�X8��%�&&Z���S0��	B<{�)�F2J�A?���a}�O\]��r��@JBK��}��|��� K�=ZF�`N�yR[+�-��V�&�!���tZEZ�A^n��Qn
f�P��FG��r�z#�I��o
��p��ځ��@q���Q/MOh�=�sun]:ߵb&3~څ�#s]R��-11'%����`y����)�k t�����T��PҤ!�WLϮ�|����.�-��&�ϯ��;*���u0/y����B��4-��>d;n�:Ѫe�HMD�~z-���������UT�� �?PMk�����9��ߺ�h}�Dh��Q`ms%9���C<���>t�^��(הD-k���]��+qN�#lG\�#[���̬�L�g���Oŕ�W�IL�*_N���'_Z�;�	ExJ(#�u�� ���Ge�xR���2�9?I��=����I����\������'o�Rj���'�}�'�}����O#E���kp�Cr81 � �ຝP�/���R���1b݀���M��꩓(�Q���jnz7�;l k莲ew����x�}q;
���A�1TJ����
@R/P��5̇�i�U�Zہ�Y���j��eQIs8�/�6����,p��	��o�$�=�oxwE�(U@#⻢mZP�0N)�ɉ*r�O���?���ؼ�#��t��ag#Q�G������_ߢ�k�
T��& �`l*v(#�+<��P*���Nn�
z�ǋ��J��yR(nNR1=*��io:p<����n���M��E�Ƃ�ƾn�A>�q+ڛ�la"l���Z���&���f��l�n".� �Z�|0�Po�l�h��kzm�nZQ���b�w��c���!d\��߳s��\-�O�L��j̾N3������ppA�.�K\��1��\�|m�c�[i���^+�.K�;��f����|�B�ޯ�3��n��N(sa�d�S^Xxd孑��$N;p�'��g�S��	\��1��h���~���_��m��ͤ��;l � ��Ux�_�d,�x���Q� ��nа�7�W�^U���=r��Ǩ�q�G`C�U�F4+J�N�3��?�ţ�j�_i��y��c� v���Y_�:�9oh�CN��m�(�{�Ϛv0;�X�����[����j���~(g��Q��%��\�+_5k��P���@��pvc�pы@�!�m��/��e mo)$�ݿ#v��%^�������hh��<��Lf�����V'_��Z���f(i(+�LI��<e=�a��u�eN�V����]r�G"<CB)r�H�〈�+ݟxP��l%o�1_�1��EX˕'�/VW��,��ූ���zP�������(�d1��76c�wi�ى)�h�>�\�Y>r�c� �-7'�"#a�6�z�uqu6�P����3wv�����F�����U�����`i����� �1Jz�	�m#�"������qk�/'��z�zk�Ro�uOQ�{JB��߷�0� ���Y���r����MA�v���zǙAZ��Ww���ytV�.�����ym��,pM�'6�f�g ��W/�Tb޶3*\�*�@���� Y#r����B�I�r�e�������0����70t�gcH$�H҇}"����,���TN0�Ԉϓ�%� ��0ȵ)Ӣ�y���������x�+aĽ<�R��Ӓ#� h���I��",MQ!	W�T���/��2�<�9�M��f��f��¾�^��x�N�O!�p�,f;��h�,��]�u�f�����:�9�E<^�]�?��F���-.5�*�'M�f`�&��vM�p��H�cس
���k�G.z7<���f*|2JI��X&��(���#�x�t�KM����Op��:HҗN�Ed���t'[p����M���il|J;16r��f��)~���Pihq��8�(��&Se�r$�J�xi��j��q��� �C��N\��rC/�Þ���-+�I�ǣ���w#�F�KRe���Ģ�,�3�0v�$��� �}�d����(bt�RA�^���;@$���I]��`���Z��ζy�_�qƧ.h�I����.+eF��~��%w�_�ﺃn1t:7+}�<���@�����-�-��YE��(�J]LcMhBg��� ����xƣݤ���0'u��7�^�Qt�-�3n���X= ��������:m�g*7��a�i��R+4[�NiH�Do_(��S�1�_����`<v�#(@��Y�-�DŤ����{�������Ss�,J������0o�	����%Ѓo`�j4p�M^#�I��<`璵������>��8�+mf�@Ef�}���#`ﮮce��b3e�e�����]�G�������wE�9�����C\ʘ����ߛ��|��z���Ȱyo��4R3��M�3���u�9!4��G($��'���6�\�g�J�Au���;p���B���˯Β<d��A� 4/���X�w]E�5��g��2����f[��y��G�f[0ETs~�N0\?}�?�5�c8}@\
;���}3�ؤ���d&Q����u��Oc��В��P�{������I���1���R�G�V��P��]˭�j1���B d�1P��b��q��<��Bm��W����\�����ĵ[��t��{�:Ŝ���i@5@����г8�/��v&P�4HlqD��\F�|��:�/��-�F�d�/�T+aq7�Bq���yīj$�RuO�y����'F����m/ 	}CCPFF	��f:��F��J!g�Z����EƔ��@��u���͔OA���v53�nA��8���n~Y���3�X����3��ǊT��/b�0Xk��,�Y��~#3�Gmw�E���
�e�H���z�e�1�H>j�43<�^����w��j�9���vT!���FN>��S� �}c�r��常|�l����}��I#�#K�����T�[�@�-}�)�0�.�2�Ȣ&{>�JZ�n#q��j0A��_�R-�/t.Q@q�ݑ8g����+����}I晈Y=���&��͗c�2c~����]�"��&4���N�vݡ�הp��:�"�����+H��@{�����՞��L<�[�nx�:������s��W��5OA\;[���85�7	����۲|!֓��a7Fu�x%i��	��4�̭^$GX4��r GI�/��;���G3u+ �?���vRu��Ę~�Y�����c����R0P��7"�##��&�B��c�hBF����_��t���y��Ƶ�@,e�2$�ϞjB�+��m��������8㱟��ޱ���i1�HF������2J����?��Ky"��̊R�M�Z�c>�'|�m:�1BW3F���a��1��̅gz�y��D������D�ֆ�s 6c�h�b�a�X����WK_n�=�V錶HSK�,�Bf�a���w�>w{Yk�}���g�̆�\e�қ;J�C�͡^�`/o��by^�u[���l��a�LM���P��G��+m�/�a���Uۑ&��7�E�kl��g��m��o��jS�\�zR/ɑ���M� ʇ�M�O�U��E�����O6��)�41�ި��8eIٶ@��X���H�?[ϴ��f����'�e����ɷa��������k�6j��f���ω���{�ֿT�8�����]n�3�VhV$v����C��%����=4���"�M��7��no���s�$Z��>�O���ފr}��|� DP�r��N?s���_y�{�;��_7��TR�W��u59xMQ��p��߮���ûH��;9�q��&}d��������A(&��[�_ӍF����Y�M��(�bV0,�I�<0�9�=k}&aA�x�]η��1[�GRc�W~v�)�Ec����3y�':�X+Qu�HD���;��ʇY�z�I���B`���߳ ���#�Y!Gk6�f�4b"z���0��qF���G�x����1�0<%:S/V}��o������V4	����D���M�q�8��V�Iz�4��r1*2z�������+ɵ<>P	
e����432F��z}-�5M��X�l�WJ5,�΀7e�Fo%>	|�������PbE�h�n�����bG��@�WEq�.Y�#�M�-M��.�]w��������g'㷿��K��k!�����џKc>u�Nw����b:�bos����xgy�M�4�������A�SQ�'Q��	�і���n�@u�89Hj�	S1V�H�nF��ȍ��NV*N�2��9���I�uO�S�Ƌ`|H�hћ���5_�ځ��Ƚr�j�;�$Λ���&#l	n:�)�����`�܃]R��!,J;
���ZGM�ۉl��.pt�+7BKg�9� ��ȇ5V�o,	��u�;v��6���_ۃ���5�-|��aK;`{8�9�&gD�s�39�z�J�C����P+����]�����1S/x$F떋�f��D�!�n���6���L����V�Jە�
�hSjc��r<7�O����xmKڬ$��}�s�U��U,����]�{o��@���|�l,�f@�iC�R�B�S> �>yHտ��@�	��w���ER���
��7�]z�ܓ���TQ�G������g�I�(��]���8�*������aAS{nS)�WLl�d��)c ���.K۪���Tw~�W����O�h�Jj檖�/�{<4�?�?���Z���n�s|��,�����U������MM�m5��^O��m���c����@MV:Y=$M��n=����Z�`N��kr$�i`}��G7N����{�"��
��A�����zn��nR����PAMH�]�C�tV�b�'�y�l*��o��B�H��:�T��3Œ�Rd|����byf�r��З|W���;��NP����]d�F����R��%�)���UH����W/�xb$B��H
�U��2�ƌ2)�c����[+v�<�Ր���`LK��-M8ٮ��V����d���C00���]��%�R�l<�m�@��:p`���e+�6A�a`�b�TB�@�l�#��5�qg5C��fS0��6��ޞ�Gbx"�:�y`[)��=��˦��p�i�������Y!���2�<8��E��G+{	� |F�;$�5޽YG��O�;��	f-�h��55��K��\�ز�$n%Lrҿf��B���+z�	��4GL�=�$i
@�����ӡ���J40���8�q՗���A�<��qI!�%I�!��m����� �M��^�@n�z]S�`�@|/����?�w��+ZC��A��V�M�}R�Z��ʻ�fb���]:WT��c�Hfa�""�wݜ�C/�m,b�i��,9A?򻰋����dj4�i}Q�-����Ub-�#�¢��:/i��󯁚u	V��7�]?�ϙO]K��J��
�,�8�y� Q��T�O(9^5k!��N�K��4MO�7�c�j�=!��J|Y��R��z�^2���e��"KYᒜc����L�����f�zq7�c�[��d& RV: �^~`�z��Ō椲�� �ŏ���.���� {�1���Cf������rH�:��><�3��ĠG���Ҽ��QHX���~�EBH`�DS����lF:��c)�|�_�\#��|���^�u�Κۋ�0��G�ČD�����D�Zi��.,��NQf5�N�x�����˳�-gOK�}�]���IS�XN�ɽ`{����L�}�|���	>���T�u��l>�郡����f�+��y���[<Vp�l�lE�T�����F���$��C�q2�dڅA]�ZXn7ǰщv�*��։U�.������D`<��O�v6Ų�x@��s!��yND��)�x�Jr�dG	�>D	��׏8w�w����Pv�H���`�������@�� ~6�E������⎛1{dyG���v�� �.�o��н�_:��f&iُ�9⼚�g�@�iJ��Vb�b���d�i]��-}�u�u��P=��/ż�P<,���Q����+l�z?��@�]Te��h1r7�0�d�6�
ŵP�LG�v�B٧M��5v>����U�
]yh�\g!�H�a:�]�ʈ����fkc�v����ϸ�L�3�4'��tm%�pei7��f去pPR��D)�ժk/�8=��t��J�51��l)�V����!≮��k�� FG���vq��°�*��~Nu�"�@��	Sw��!l1� W(	βXQ6[��M> �m^j(�y��N�d��*Q�͡�/��d�a��8�҆��! ��Fv��I���)X�Rv��A�qϵ{��Q��@Bnwy���,(�9��Ԃ�i�k�أ�INsb%���A(�.V��웁,J���=ήN�4M�`�H��/ O�f�>Wi�~����&�oE�S=�BX^�OKk�s"EK�c��n�C<	�ގ��ۥ����2RI��mF�n��~���|''�&2��c�am�	)����8�~K�4OYp2T]�/C���*��,V�u�2���Q% o%�2�������f��֝�P�C���LM�q���0�(�b0��?�ZT��i���\Mb���7�l�hdw$�lHu��5=��6��������H�ħ����0��O =]>&*�_f���i� H�c6��O����u�_�t�/S"B� ���훿c����f��Bo�ҭi�ap��a򐘀��?9G4�W�'���$�p��ԉc�KPF��}�:�d��r��t�wAÌ*�M�c�TY-���5�[�MH����ǍΎϐ��!��As���#-�>���q��Y��d�\��h����� ���\p$h�Q���>JEP�%�`�*�G1i6�j�U��*���$2`����qÝk^�˳5*�a�Ġk��Df�0W43)O���C�ſ�����v��D_T��t='gM����^K��"C�G��4��i�2&*~�C7֢D+�n�:c���qPFC�Qlw������
�ܒx����͞U�m�|���}H�5d�R2��	3�VY9h��<Y�Ω�(���@�]Qy�-PN�P2��V�.b��xȔt}+i���Q��{$�{��O��Ϡ�A(BѨz8�ٯ�tH.��<Q8�6n�D�`�.�BXs;�Lw�����n�Stg �w�����^\-�i�������&J|���y�׾>�3��
*'���� �f�HER-M�b��r���RF~ύ 8|D�U3yI�c5�A
�:3ZG퐈F��Z��������(��{�Ǯձ�KkX����9z~@�"R#	�g*(�,E�Ə�y����o�&;S�+)�x�b�
Ģ�8ͤ�@��&���8��k3�:���{y�[�w�$�}-�������,g�D��Щ{�sMǞ[n��4��&b[�N$��uT^�ڇ�k|��j�Q�Y&{�l��V���R�u�T��Sڐ�SP���]<�ݠ%�\am�����M�(R�b����h���!mX�Dꢠ溷`{��0�͆_�ǭ<�H���V�T������hHC�����ݠc�]OWXQq�X��4�xU�L�5���p8��s��!�%2�T�Ҍ�C�]���>���0
7jA	����v��S������I�N���k�Y��Z�P����t8n�կ�/���u
uZ����Aܚ濨�N�[R��{N=�0h%�@ذ��J��*ʕa�\���������6a<�g�8�˪3GS��iQj|�����|�����
�2(�":�hl�~P��2��=���R��>�l��i!��\R�+�P{	^�:�@�0X�\`�=S*��@��:��M^�H���<CjЛ��F��HJp�
���~��خ�P�s��EΉ[��#�ڤ�S��2d@�K"c���n�5���*�p��<�H��`i�vX1�3���{�v9n�bn�E��e���Bg�D�<�w�ʋL��5ԣ����3��:�M��d�9��0u��,�+{:�����{DSRi�b�a�����9�IB�ה7_��+�,�ԔW[Y/���H�����G�C?5��+�άsd*�@�.��~�
Kʃ�o�?�YV>%`b�OU:rt��/sL����8B$��I�}��������l��>�3�I� 
�U���NN%�%L�	C�-h�%����ʻ\S��E��k�(�k2[?����7�; �NҊ���.��v�~x���d���o8�M��*����j�k����l5ӝ�q���\k(���	��J>)N��`J�[n|Z����L8=] ��pc('��t������v��g(��Bb�M��e4?2���[�óہ��Y̮뻗��Ⱦ����%��l�wx3g��ߣ����w� �����^�˽bC��{��t�?���������W0>�W���t��e<MX��CAHC�	��[ڎ��Pf]�<��<w5�a��:�
5�o<yQB�5;T[�:ܗx_��f�
�
E�s�}�aGA��}���0'e�!؜P�c��s�V2cCr��-�N�|&�J������jY��֓�a �R (�r���i����jm�z�	 S�z�|��&�W��=�P��cxɄܜ�W�a������儂�|�|�P��	\+�˿�PY���I8��rۊ��X��J����Q��@�2��=/�KZ�>�v&�V����/l�b0�iBTҏ�*do��~�g����]���F�^OZ�w��h��������ͧ!���GGߗ�����鮸$A��r�p�jU?��'�!����{����G��>}��
m�1_����g�'�ŝ=� �ؙ![	�X#���t��X���y�oH˳�RxjRi ��O���xYه`�1��b��3���b�k�&���w�ŀt��$���w��N�A�o��)4/~mqgr(��c�g�t�Ϩ��wބ\b
�7y���U����gV?�&�rKF�XJ�G�VZ�}��r���v1]:��0�f��t?�%����,������-2dFz1�3� �վm��+�T�u}�euV�Fhފb�{��<�;�W���&;�㠼�v������y�����D����DG[����9��U��	�J�hqJq�b�?�9M0�,�+����i����)h��Q������0s��:��9V�aK�7���K��-�R7��)}ד�����c��w8О��rf��[��qQxFG��_Q��CS/�1I���6��C!�q��Da��̗e�p)f�+X�������H��2ʳgǑ�,�%��D��l3r]�,�tw�b�.�����\K�����Z�ԭ݉��,��؝��ʃ'LAY���^��7�P�|Q������lZS��f�� ���e��sQ�>l��DY��hغ���2HV
県�˼`���:5�YW�j���ѠRd�l�y�r@C� �!��n�R�*Ϡ^��0��>��;)�>i������o\.��Q%�qBxa�4����7��f�w�*"���j,[�	"�j����1������RZ��L�d��:�����JWwǧ� ����+���|�1�|�$Gf�8I�&H�P�cT�,4T�Q�J�ެ����v{'i�ʝ�a��C�%bU/��p��6�V�[�VQI��P�&��we[�j�K�	Is�,\fxK:>����_�}���"��čI�~��Q~蟳�z7���њϬ6�A"��3x�x���\�:�0�F ȿ�< �nc�-;kP�Es�ݯğwZ�'L�}�4�������ӡ�1�T�JD(˵ }�G�3]�iL����Ȧvj/�@������4��@Į�\��챻xV���s}�R��h�vS	��v�
�����j��̛S��~�H�6�{_�E���JfDIO� /�������ch5�	�G�%F�� �Ԏ3�jKc#�A&s�����)Z�]⇄vg����g��_��%��zJ,�,%�A�;ѹJ�) �Yt&ww�`:L��V�{���S���3�d�k��u&�ϸ?�@R\�\P��*����g��k������V��g��J�㫝67��Z�W���(]fYi�p���猴�zLR5�����1�d&v�}�0�z����b��Սو�	^��ֽ]����$��I}	�����>-����d+^�7Pu �2i_���X6g�6�D;��ۮ[[�$����5�����2���*���R1Z��r������}��Sz�N����;ޝg�����]��v�?#a3"�s�i$eD~{��>��q��t�%j����SH��FѾ��/;��S�v����[��H�i�+��c/�>���![�˸�ɧa�h�u��[�m-<�b)1dB挡{l���"+=3����/EO)4��6����>ԗG��%a�el�Ѱ4�]aF���j�EPy����%
����#��p=KU��8�ar�B̩� �T��=�?B�I�9�+(i9�Kq��'@Mw�F��@ڊ{G�@��%Ђ�8M�}w5h�٢m�I&���9�?�k��ղ�`<����`xB�_��O7�aF�<�;.A;�j�CK�i�陦_�{��@T����W�	t:���� +��G�#�/&��,��*m�Ffb��a/����Q�����` �����#4�����3��̊;��h��W��q"(;3���ρ��������G��_�{�6�E���~��H�	�S'�m�*��p�PZtV��D:�+�Ǻ64.���s�6%P��^[��=Չ)s\��o}��� R���x
�S̻�+om�k��FBF�7᮷�2���1��9�����X���>���l�֘ǫ�G�:X9՞i+,l�u�b:zs=.1��|� n�/���!�!�l�L�KO�[�œ5�A=6u$L��&U�R�8�nd��&� �~V��u n��5�\#�ڎ�q�
!*w����v��L\a�U� ������.`��?8�4�ӳJq�g+ÿ�O?O~g}����h�:��3
>1l�ߦ(�;�09�w����x,K��?Y��݄&F���F��z��)*w;R*��{��į���x�(�z�m�H�2����wY��:��9%�I���*����y`{��Q=V�S�1��X��	��)%��iqD9A2E�0q�+�[�LJ鿨�3�}�]ݼ����wb.̵h4���5�$V
	�����­�H�D
/ �zPP���W�L�p��
��Oբ�:y��j�u��ϑ"F�G��1-M�m�I��e��*l�?7��Xh����E>��(T��u`�j�R�}�/��LP}� ���tU���#W	�En;�1�Θ�+���?�U�G�g{kW�q�,�w��V��f�֏c�^Z��m��h��M�����E��X,Z�����ި��,M��P�>��?��48�-����4��rn���*\��ɽ�S�:7�1g�N�Z�3J�� f��>-�8��`�-Ҝ��\�F��Z-]�JTN$�l���_�ǥj*Npֽ�8<cPp�k�������pS�A9�_��� dƻ����*'�\mo9k�c`�`z�H"�{��J����?<�=��fs�~�zw�o~��Ěp�_����"�T��$�i҄��@>?�7+HӐ�����ɾ���Mo_eb���=^���Z!�,���c�GRx���k��Ւ��uM�Aҧ�G��x��;�
ן��i�t_������\��h�$�T"��/����1�i��N:��;{��s�{4���,�ik�ٗJ����%���{b��_=�Ny\K6~�{ޔ��'6W�|��,��U�F�
Z<�ikdP Z*����Q��t��# 3�w�1������x�zu�pu���b�Aлa�2x���9(p��7�&�'���x�k=p�*>��?���U�AA�� -�c��V�F>aP�#�����:Ȋ�U�@�����-m� y�+�Z��<LVU�(�`�F�-XQs����U��U@bOD�x��]��d��--⛗LV�o�(��W8�s���%Z�X;��	dZECWzÖx�`�]V�20�h"p�X���=;ƙ���4}�:B�$�*�����C|��ǧ)�iy� ����d68v��:d�&��iu�zf>�L�C�C_6�-8d8 ��n�%�
T���%-g�͗�ٙ�����~�i��)I_��za��qS	�;b��>!�J�2�W[�MގU��m��c����Ҿ���hC�>	�M*�Z6� w�����I���YX�Хdŕ��n{8�:EUw D0���M�&!&�)�@�x���}�f�w#b�Ӧ�U��i����?XI������pZ��:���O�R������ث�k��&~�"\"oʴ��P�bg�ʐ���݅v}*�V �"\X�)
���p��'
\|2�Ũ��`��	|X�)Gſ��k�|]���ȸ֔@p�*}�_����NʠR�M�T@�g1�@ΓP���B�/�o�/��+�`��U��`ݧB�k!�gu��Y�ITs�s�8M��_B�vP<<�!�o3��m�@�ι��O�\�@x�$Bf�"ç`�k>��	��1��4�\�R'�NFA����]�3=�������d���2j�C��5Û7��֮�B���ѽ]����BS��Y����4,��L��+u9��J����
��E�ph@�6��Ր+Y��t��<H���8J���.	`���B-\p��XJ���¸
����/�C��'N�r�Jv��BA����%�Z��K.q���`&�6F.1$���j�ď_��x��yP�	A�C��Jp��J&9�2�\��>��+gl[�\_s*S{�~�e����ak�Ɂ&"F�Y�1ø�T�|�E;@�H�@�T�`W0:�,���{��
]B�Q�ޫiW���D�,�R�D����R��M�B)��u�ez����<���FJ���mM�# �(�}P�6�,�Tj˛>[�Q�ƀ�t�JKV]1�B�l�����'��<[||q�� 0���h�A�qV�����K�]�yш9���z�=>�m�tUHK����F���,�8��}q�����>n��E�h�ʀ��Y�a����9v��:)P�K\:��,�Q�N�{�{�U�AN@3DM�/����α��?x�m�q��g������r�ݣ��t��h�Zn�q��=ٝͅ� A�� �ѫq�'U�q�^�'S��-��`'��]�Q
�'�NJ#?�v���3�F��"��5�S�p���]&��<Ϟ�)o�Uv�5���{rSM4i/zT��$9��TN'��-�.�cu�ҶÞ�Q����q��.��|��:P�:?i�����V%ɫ2$��Ǯ(D�k{�z��rƭ�
v(WS��zf�2��;��̮�j�A,�qm�5SS��Af6CWvb����ب]��8���y���i�ְP�����hr^G�>�!����ƪx��N[�ya_�M2OS���Y��i���B�^}g��x�c��>�LDȟ�&?�u����)���u�RĐ$%m�Ύ����k��ކ� ��1� ���7Z����;�]{����@7.�]m�d
�?{#�"}���"�����N�f?棷C�`�`co��E�g�8ۜe��%�5 Q`��� U�b� ��e�'�v����`۾[�G׭z�}/�_�c~|ܑn��C���x���2n����Ľҷ����D��͈��+.���������g5���no5_%�;��4y�?���<��<�U������L dò!J�4'?A�Tzz�*/BI��Ջ��`>u��X���NZ)XQ�.�+fJ���oS��._,g�� ��u.�0�P�]�U�_E��A��w�8���M"Au� ��u��}+��yg�V���Ox\2jqi�x�|��ՙ`_�isz�P�&�#�'�D=! S��NѴ���t�	�s���D��0��Кݝ<�A�6���uo|��wa�����C�9#!SȦF��n��_�E�����ױ��0�&��JpPoLM���I�!N�^���[��t9�C�;n�!�i �3G���}j3��}.�|y�o�,�Lzą��l�u��<:���= P \���8Y�f���DP�(��}�-ݣ�q��n�%KX�uU3�Nh�W�����+��[���C��of�d"���@3���0I���ő��]e��΄��)�����k8�F�@i*�7�ћ]�俶�b�Hh/�z��g�o.R�5�]���%�	�C��h��@lk�f1��&?�4L�&	y�b�r������M���i��l�����
�,�?�&� �P���������0{��5ru���:3��k|'OS���⡤�F0�r�D�D����D��f|����EC~�3�|�Ç�<|5BW5	���-�[I�)�l�!�@��`��s�����t���.m����;h��G� y��2��G>w�%�&߮И�%�A@�^!�u���,g�">��A�y���=�A�:���d�1P��^���q`b�����삃o^j���*K�w��7��Ne�_HC���O�]��ʄ�Q~fuL��p�@�gXv��@]�{k���t���b3�=U��Oe�3�*��R���xj(����g'k�i71>+�-}�"ϙ��6ʹ�{չ�ޟ���}��ȱ�F������uW�1{��r(h����uiI�y� M����s��b獼��,� �h`e� ��Տ&��ȭsi�Y��ؐ�GIQ�xժ�`��0�Ɓ�I��}��7j����à��WP��_#ۏhE��x�Z�{��V�ַp"LZ�{��鹦R�}о��<P�ǳ�/��@����!v�*�K{/1w
�	���?�x�TwL�}fǭ͆�<w�(+e�Z��-g&`�-޲U9���>�M�+h�����m�y}�|��T�y�m�}6h�?�"��U�?�Cl���J�3$]&$�'וy����Y �Ýn�K�L��u�F1l��CǛ�&���]��������ʡ���ڞvƞ�k���8�=��SUvL���I�&S[�����d�?�n�xz�T�?-f�6׊��]Fb� ����םQCݐW�_�c�U��#݌=x��lqah�x��Q�����y�\BF���Fk�PP$�R��S��XO�_��cb���s$O����sN��:�{|�K�D
č�ҙ�ՙ-P��
,�g(��Cb^���ґ
7*��u@���7�t��+�/�Q{�j�������*���Է���a�ѹ��n��Z�U]�1�mEǧH6�R M��&���Y���gg�E��+C�}^�M2d~��3�cP�m��z���e����N���������WB2/�@���U/c��K�1�lx+�N'�;��~�wl!��ǻ�V]�N|;P�fg�w���Hf��Ül���o�_�nCx`���X�7 {� ��O����1䐪5��\5jD����������D�F���s��Mzx�1]�ثX̎p�0�׷��5����^��� V���N�.�������!����d��[ʯJ+���^����*�hMEm�F������ӞTn3l�0��흅��-ed�VҺ�U�F�m�wusJ�L�_4,�
�P(��b)��;ዟy���<�ƃ�.��'�- N�eߞ�>,�D<���%�UDON��+��ؼ̆�R�	��Bތ���<��m����"��'*�Zh�� t�IM��[�|����Z�.�ݡC��>���M-w�!�ʥ�׮ڐ��*�*r�����%e,�D�?�б�m������ۃ;$j3͝�bq�51��,Ƨ71J��U�`n��O��al�I�E�VD9sag�Y���>Y*+�ϕ�a�C��~�Q��}��a�9ǻ��c*Щ�L����mP�j����V��\1�e�-k�9��&�u�uAfB�b�J,$o�^�%~Y|�R��:�M����{p	x3Z���es������x{5;	]�(TT�rv9|�b��$�<�1m.���b��㖫�G׉�Bq_4F#q��2\&Қ�A��v����zmȢ��zp�.�-�^���<[Sܹ�M�v�(�v� m�) CU���,�̱�5<I�S�x� ��d)51�@!C )u�.�� �oѤӈ�t�j����Cx��+P�Tݮ�0��R���.J��Z>I3W�f�a#w�D6k?Q��J�)�y�fA�@�!5�]��*���߁�3i��ܔ���n��d���^r$��6��v�����=�23T4�w�*Ey��ZJ``�$�)�q��gB�c�+���k��y�˅������Z~D������X���p/I 1������t�rH����d̂�k��'X\>BΔƌr"����ՠ+p���Ua����a1)Y۲��hB�7���"o�-4 /�|!x��7�-�+�K��Yyd��j�«�o� 0J�?���
���m����Y���+�i���ך���FZ���wgr҇x.��y��������209����Znͪ�C��c�w9�F=��1\�i��Tt
������m��0Ka�x@ �ci	�Nǫ�P��,6���8y^=�P� +��+�[�E� +D�.=F�x�u~��rH5�aqp��8�gS��D�
���:V!*���:�#�R6���+y���L�$�V�09�9���%��nH�N��O��Ķsn�yZ��e���<���,Ъ����G�t~��k۴�X)4�آ�bM6��U׷��������( ��,7�X3!��~��NZ�+�1'!ɗ�3��Emn�d�IC#M�j %��2��_�!&�~��Q~x��$�����ȣ	]0���	�B���M�A�����m��Q���fW�� S昿����~E���|;�C)���>-���.��c7=����vØ�qN����f�IL�,�g����E��׸,�R��L�q}�2������Ek�S����������V�x�^е�h����]��D�j�}̒�1Om2z+�e-��4�n���Ҍ�r���5��r����G���E6`������)����u�#�Ӏ�֌�C݁}I�6���vpV�n?"��p@�6���x芦��΋^N�;,p��q�Jdv��*bxZ��+�]�F��o��e?��V�-:Sq��%}vM��*�b��'n}S��.������z�X�Z�6k��7��tܜ.����'��C�K$q�T����q����v�J�-�(��F��zI�?��&��0��n��L�#@ ��\���8����op�,4�[*�G��SN�,��ČU�C�t��_������ׅ�)%�z���S�3�;O�'��-N����U��f�m�#]��a�GY�ĥ��yK
�y��@ML�����Bm�  �6^������nV}�ב�ǒ8^���CC#�v蒚mn	���m���D䟴��B���^��0Y�X_p��Vy��j����W<�e9lO�p2�e�c�Q`)��c"�^̳=9�\�`��"i+<7�C��Yqr�&�Bx�.��.���)����8L˓eu8N]z�7�k�3��2z?P��΋�<�]��U��8�>wP�ZC&0�fc�\~n�)�.߉QD�i\^����\|(��
�-.qU����Z�/�L��>k���}�-�̾g��?);��\�*:K+���AY�����Sm���)g1{.y��r_%�6ӹ��Kc��ﭏs�#��2���g"��@Ӽ�
��A�T!���jͼ3�
j"S�*u�y3v �l@!0��~c��ȅ��^n��[c�Ĺ/����n�5W�T�W�n�˨w�?Nv����RO���,fƿ:2��ڱ��%�����J�W�#��ؖt�|
r �61X+����^2�4����[/�}�6����hXB!y�|��x�N���<|�$�@#���W�6.öW�E,�s	>�x�-￸�nM�s��=����;�
^����bX�M�;ԏ�3��X�T͙X?��͙�w�����o�׷���
7�4�3�G�����?�U��W��	��v(B�~2��іA�;��8�m�i
[�T5NCZ�,�Я�уcF��I����Q�=��_~��U<�����(�� �.����ﰊi������WMq.��T�i�Y����L��RO`���-�*-|��y�Th��H�p�i�����q\��i��v��4�{wZ�a�
xk�yDV��n��Y�P��}˗���5�O>p|I�Y�Uӻ�X,'GØ�W��>��T �L�鬅V�Z�F���Q�	k:`���=�H�|@��A�o�P�Gk�#I ܬ��NlaV�Ј�/-�e,@�PSp�o�Ѕy�Z8Lؑj�C֏�λ�8/��SK��,�fl5vR�XK��7�6z�4��ɸ)`o���v2�!6�/f�p>�Nrp�m��77F2�,G�_p�*�����S=u�/��y�8śq .�$im[�"�&zͬy��mIb��kWY���(�@��P!㹚�tZI��ôY�9ED.���6G\f֮�jBC�~�#k���IM"&_+=}�P��� a���YPL_I8n�#���������+ۥҷf����G�d���Į; ,��N�H��G�[`���yϪq��1��/�� ��I	����eKr^��u껥%,`Ɏ~�7�UA@Ԇ]���HxL��r"q��������e,��P9��R˺K��PJ���5�W�^he{�g���/����nړXYfE�?�>���J"�\VU�����u]�-JbRZ˽�)�'G?�>
Ŝ7��n�p|�̥%�����4��1Yw6��:��#>�E0Xqe� b���جݏߝ�Գ��1�D����b|o�+A��๧@����җ��8�E����51W�͞�#���9�L#n3+�;���2*d��g��A���c���o�wƦ��;����0y+��N?���Ⱦ�(q����8���M�I���9c��+W�|S��C�����{f�Q�'#�PJ��)�%���NW3�^�b���_��$.�s�ж�^ߨh�a'�Q]�v��)�'ؖ����7JXw	��0��9]p��i�M8��� H�$�3ѯ-�s
jwc���h���������9������-s��8���u�B�]��+��U>������7�~�T�{�����a^)_b�?=��Qm��c�����᭔*u��r�T��$FG��ٚE&g�]�rI^��3N����C^�[�?pҞAB�mF��nx3��Y:"wl���=��������t*�dVQg1.(>�n��np��`��Ie�L��9�w����I��VKڦ\���� �ʆ����͝���ԛ��A2��[�j���[�I�G�0�m8�$�8�5�Ӯ�z�6��d�ǋ�ƺ��� �'-=,��D�|?���	��2y�V��P6�+��� #�p������E}�6��$�����`�ڢ�ᐓ5lN��p)�+��ZFF-�_�7G�_�"�XB� �z]Gx\��ds\�q�b6 H.;eN�I��/�Ƌ��
o�cPT7��wg���e�����W���_z{Z��X�I�CL������!����{���y���pd��b��7�#+E������0���pɣA�����: o\=OP����A����[�0�ǂ�F�U�O S��FȳIr��ZA���:d��HR���V����u��+�Y���Yv{�|�t�,�~�Ce�"J�+{�,��F���<@z`�U�?��~)[�:)p�-�~�^�+~*����q2(~�f�Ɲ9�����ӭ|���0�6 �rY}�W�X/�ώ�外${�w���dgZ|����.z�h�na��Eʼޡ4�#3�Sx}���<ɾJ&#��\6.�1���կۏ@0ϭ�񭩄�`H��s�I�3� ;t�C�I��v^�]/b��2�;+/\r:K�hA���!��Fq�E	�}�$�tR�]�:wM��Ybz�e�/�1Jz!3�����@��H�NJSXf͍z`�nV�	v,�F��&��_pQ����G�v���b)���Ş�@M����gf���m ����5���z��%D���q�[h�d�*I곩�X73\y�G���o��%x�@.�!6?����{ׁz�=�Sw�!��R\Rï�7��t:���UJ% ���E꩑[>�+k@T>�D����N��-Ęz�F�WY�-@�%'r9����Z���t�(_�u�</��t��Y\�I��TXK�9aW�Hd�G>��a���?}nv��_�Db3H�"7B�5���b[b1���3čc�{J��-�����m�l*5�ω�Jn4<]�+��o��+L��	(�N��d}r��6�Ŏ�g-�04S`SM��a���=�F�Ī���(�����h��o�,}���R�Q�
��߿X�o�r�%Ǥ��l�>�� o�$V�jX��;����+r9�%�����q����\��m��A}:�.�$K��0�#{_�4w��
���MN�H_.�p0��"{�"5��>}�h��E�9{A��Y["~&�;������ӈ]]�dl.G�<)�O��T�d���tb�S��I	�	��F5�&�C�b�"�;��^�V��C�;v��)��]��u,��[7�;�#�鿵u���z�6����s����.�U�4���JI�F.�w�
���%-��GBn�c�[����a��
��7��21�ꪗs�0�!�Z� ������-�18���?���򉖟�݌�P�
9���$� ����~���l�����H�R��|28�OT9�����b��i�$�7ٸ
7dJ-�6���_"2!2��R�3hn�ƃ�Cx��Y�`ą�hH2�B�����b�$��Jw�+�zR&��r*}�	q�R(O�Sl{�J��Ra��k��ck�Ť�X�q6 �M��~��W^Ԏ鷉O�$Jǵ����V���@�����!Z�>�HV4�:X�]�s�8�C,�^G��@��w�Jt���[��_�@wIh��ãT�H&�d�J#{�I;�?�'~ޡ�E~T�eDK� ˒��3�Ͼ���{%㓺ӻ�p�?2�� �S>�Q=0�+&�>'�0�ZO	W8��T�ss�[�Q��Ա��`	]���������}ނ*rd{��a'�N��p?f.�T$�fY���8uB��0RJ+��ދy�$@�8�ի��� E�#���������cڑx�j{�X��/p\EY�Ψf���\�h�E��|�	e7�%-Rf��d]�lĕ��GM�`���Й���B,�c�^��xI�UD�r)Z�'@�b�gTU�	�� ز����C��~�l�� 19}��;�����˥�d�ݮ�3׮��ɼW9z�.����pL��*�1 �"1������� +G�U9��'�_�8K�0��7	�Q�:�;fA�z4٠$�k��U���F�LOs+�������9��J�G��䅆˿2�KSAS�k����y_|����T,x%Ҍov�P>n�/��X�`����<����	����Z���S��Aq��?3|�����/�;g���Y��,3!�_�!&���N�
��ߘ�4R�K!��K�v��g�l�����������cr��`��C|���e�/�b���Ij���+/�5���~��w-j��k'8�NP��B^~�`x�P=;bd:të������ә�&_˹B�,���!jk|3���q�i�x̛�x+)(�"ӖbI���l4'"�� 2�/9��vK��[8$D����:�T*�)f���	|��t�FaP%]C�y���.����3m����yܐ!��[4�i��N�I�ॏ+��x�[���93�5�?�K���������'+�rͼ�9���\�}f���n���3���)�B�J������5��a���rŧ�OSE改��#�[��O��NճX�r��H�k�(�>��#�rTA_�p4WO��(�Gŵ��8�F6�5ɖ5����5U�NY�����^c�p���BRL1�4AE<>�*��ן��Z/pYA�6��k}�
�X����o��6�c)׽@���7��Ґ��s-�;�������)�~ ��Z\<�K��[Q�l�lLp`9��#�H�`qCe�ћ7 �	w٩��]��H#��b�9�ɗF2�U�try7��z6��ՑF����� �㲉���uH�4+"���o�1���cAlWW�Oga��5٦#�E�L�K�n�M��|V��U�+�"6s��Y�*}Qw/^�	2�:�r	P���pq��jļh�˹M�����B�4�s��DW�q��[l�?�q�� 2D뀵�^�����B."�O�܋�oe���A1����i�Zs��
12���R�W��2f�u?O��c(dk�8�u��Z��R�_��\��w^�)�9,��-�ę@����|m5Y���)��9���ƀ��2�⩵M#�Ĥ��RVC��N��V�������"��ƇD���۳���B�����UOQ.嗿�.�A��P�-8�8@�i�G�
�Vc�ىֲ��1���������ȏ�m@��@����C�R��&��e�����i���Z)B5[@j9�ܸ-> �]���W�QS�<�~��;�4����Lċ�Ac����aBB�oN�\p�nA���u�T�a��BX��j�D�>��ˇ=l�d!zTNP ��h���-nc
t���I pGܺ&� ]�	��u��ٛ2���$HÀp~S=݂68��MY��zl#y�J�,o=�2/�~�fr���;E�^���pa�D5dac���I�!m	?��gý��rK��=���y���iO.�؋zօ7��)2Q2�+��l(�;:��������SXh��������lH��Q��s��zX
̸�"�]�V��t�@�؉�����|RLĒ���ۡ4���Y�
��fe���&r�C2f��kZv���!�����w�0Y�4s��Gm4؂�)0����~�/�����0̬����l�<߂�M0G"6�D��S{��_˥����S�Z��@L/�-�o�-�˕����<d^!�u��єM��ٶƓ����F���W�)Ɯ'�1nE�\P\�2;��e��xw�PoC$�Ei<o�Y�*ʙ.@���ȹvƂ���pk����t��@-�S�(Q�����9Iu؀��$1�X�&�%�����_�$���%=.2S��Q�꜓'������ജ�/�	z�kqjØ�PN�YT��@��3j����*ś���µ ����w`�@�"� �:����J�slcӁS<~�[�q5�:#7sb�V���q��d��;^�)5c�*�>�+H3ҋ�h��W3K5��,ӯO$�Ԫ|�&��T 8\X�&��Yk��
�P]��w�PT�n+��q�h����6�vk}Y����d��0η��}^K�WO��t��5N � �9G����̤6�k��[�-y�H6��eH�.cIE��U�G���I)+��
�a�
H�U�oh�%0{����B���(�O����4z�t��)}M�\��8���R4!��e9��$Q��7�)JNc[��9�%h-�ݿ�Y!}�
��V{�$���N}\ڹ�-�#�WSc*`Lݴ�NAm��ݎ����w �ͪh��\���h�V��(�RzM��z�\�����2����@�.ݰG�s�����oV��}��lh����{��6v��������s�N���gK�������M3zd����9"k��t��DS��L_�uߎet`���)��$W�L��f�qMӄ���ԧ̠l��*��p�[�t�'�� �"쪉3��r��<�z���Y�`�ն��t�fK�Y�_%v���&���@�]��;��s�������dqm22�^e3�O�x&r�Ed��1������6�ۨ��K�AM#�_J�f�̂<]�R��1�e��.�Xl���ه`R�L�	��Mȉ^b����/�O�H�+F�U���u9+�)��w.!�\Ba����W�Tg��?��R�M���� Tܸ�ǖ/n{(���r�s+L3:1j"ׯ+b�1k����`�koˣ#�pC���l���{e�l�Li�>���zW����_��F��I4�whP<j��/�$h3�-X�U~��-�T>�xP9ླ��S2��e{�\�����:��w�ƛ�`M�ac�d9o#�����Zf/�C��C�a���l�'� �۽�\k� G+�\����l3.�Ȕ�f��� ��o�W��7ޏ  g�!�Fa��',�Jn�|��	�1 �����ԺA�6����$㏄f7�}���PD�$�zq|�g �Aꖲ́��gB @OVk�(*�5&�P���ͷ���Rk�H���WU�󉁎���D=9ed���P�]��g�y��������p�_�7�Ѵf�Z�tz�p�]�jUD�Z��5�{w�v�<��I�!-��'�b�y�j�:�/a���~�� }Z
��j�-�g3�!u2�����{�$�ɈmX�㯣 ;/Ypw���"fr֍�hF�4އ�`�ﰫT;��&�������ʹ�����P+��U�ś��1��_��������Ul|�&�r�8�����=��p6EǰF���u.Em�����P@ ں�����w8�)�V��1��Ϻ�F�k�[�,��N�K\����j�*��9>`	�4�- �$ S�Pر���='/�)8�FЮ�?�O�n���������n������]ǳ���<)"!�,=W����8�U�\�.\Cp�U{��{�	U���Lm3�q�<��v��ڼ�y|��ӆ���
��.D��nbeQ�k�6K�x��!K׾�r^����JCf�G�e.�Я8(�IBP?��ow���H�嫌&H���]�v�V�\�)�!��UDj�co<A�|�M��qE�u��zGo}!$-�?��0�L���,B���]���N'~�f޽k��p��*�fv#�i�_N����=18*���Q�.Q�{�k�hr�/N5o�@<"eL(�[�r|����4oV����wb$�wp�wP'�h�.���J �qzYF=�l� ʥ~7�ƀ���\~v3�6��a<���Vb|��2��@��D�<��`�LS�3};%�bD��D}?�a+�(Ӌ���P�b���^�֦��DC���J����f]�|�h����^6�1ª�OCв)%�G������%k��ùs@?��{�ͼ�3Y�V:�]<�$�VŦ0h��Ҭ���J��+������/�ī؍d5�4�#>RΚ7�ȍ[72�w�v�]p�;9z�	�c6�[@`�՝��w�׀=CQ����{<k'�(|G�TiӞ���*Y/�$��F@T&=R����"�z��t�ǴJ����L�:O�Uj�+�AX����!�jŴ��M	ç�xC�Zʤ�0h�x�K`�pܒ�`(d96���m��vx���$�������c>�]��;d�Y;+%\��0�������x�.��X��m`m�`�*~�Ќ�nwA��V�P����\�)rf�$2*�R8�\�,�aZ���Ұ������經�8�7��?Ύ��0������*t^����6V'Y���<8m'D�X�uH��c���� }|��	S3������n�|k$�4����� ��>F��>��Ԁ���:S��{�+9���8t&8���p�B�Y�/^}�J��L ��L��Fʣe@n����d�G�,��r�av�jd�B��0���q�(�@G��i����R����e�qP�aI�	ON�ˎ�:Ȇ"K���q��ل��������I���0@�?'�Z��&���y�)5��[�B3�?i8N6�):�SYP�»7$�� j ����t�V�DQ]>L�q�pk�*5�	�`[��Qw�4��zϢ�>���_�U%.������=�6Y�	�ڏ&��h�n?�B�2|�-������_�t�Hoʟ+@����\'Q���__4	��\��)'���%p����gx���-QO=is�]�D������B �m�dAZ�t�x���(�E+��u�	�cGB��P\��O�\T��M��3S��Δ�v�G�^�1�K��^Aq2��{���S4�6��Q괻c��؛B���V�g6��5]зq�<�������;��eFgʳE`1�U{�ȅ�q'5ܔ7���.
-)����&Ymq�P�W���򳤉Y;ʠ���f���!`�Ìv�(ٗ�{��뀡b��;Cx�[L�5�͌�rKsߖ�z�9l��HB!��:�
���Kb��5���ץ��fQ1X�l�A�g�8k�/�v��(��RS��̲������w�pk���z@4���%$g�	�M1�g�$�(�2�������"��n#,�}��RDD���}'�
=�roST�K�fH)ғbO���2����u�=���va�w��.%��-Q���6���0m�uün�û��X���Wڢ|��1�?���zg�kJ��5�`���>WAĜ���	��?7���mt���:9��h^i���N\���o�M���@�о��MH���n�}K35?�v��O�4���i!J�g�\k��ѯ+�(v�#��Dq�Na�	l-��*��_�o�����b����
o�|�QZ,5�򗲺[��W]w���};��[�b)Ѵ�b�͞L"����A^Jԡ��H�[�Z��I
����#[%��F�ސe�U��!u$ Mq�+���v�
��Rv]>�kڧ���`�O����(�-�θ`�`�<��M
��}���7�v��`!�a%�LT�c��5���Fgp1�\�0^&�I{'���^�#�����c��ha��	���Q�t�Ժ��]�Ʀ��:�^��P��q�ٔl�BSМ"�ڬ1���'�x���_j�K2�t���']h/�hJ|�G��!
|�Uc��ZwMc��	,�`V�`\�b���K���LF�����*�)�{R��ڳ�1�O��+�qB����gr�����-���~����l�ĸ�P.�������H�s��݌�R��3�.���)���8'�R8��垰S5��jYKI�d�H�M���T\��^�;17k$4�x�Ɠ�a�9���y�v�\r[�Etנ�b2)8ڇ'0_�t��ۖ���v�ۙ��bd�Ǐ���}�| 6p��K�B(Mf�Rb�u���C��s�I�Nw��X�{FvKԑ�l�[�`�O^&��a r�dbGFy�n��Z�&�_����+d���I|o��}�>Q�  @ץl�)u8T�!c�E�S����^���]��fS��.-��D\k�2�7��\6<\\ccx�<	��8�;���^��7g��?tY��l����n��\*v��up%����Io�5v]��wWmg��y�,���ٵ����z4�`���OP�ƺ�ti�no��UUTߴ�
��<�Δ�DiQ�~���Cp=�7$���3Ufb��,_���ԓ��˽�D@]���MAp
$*9�����N�G׷]I�!���Fєf{��cUAY�Mp���'�A�"�����5H�J���.t��f����|�;�p%��a�{B֓^S�%�|�}�!�켶�~��"�	G�C*�&@v[)������TN��XcV���;��C|�]��9�O����=�R�H���`}w��Y��R/U�yu.��`�ѹ������~���+�<�pq]��H�8|���ۻ��)}N>��;�h�T����hB`g��ծ��Q��s$���y��\�yc�-�t7�ok�@�"��b��"Fp�@)�IKdT˒����(��Y��'��y��#�Zi�Qj$�)���f�*������>+�i����x�����pHdz{�=$���M���F��}7л�ȡ��d~���f� pw�p�z0P��`�S�ܷ��������p߃���s�)Qu�G����kY����YC���ccĢ���w���w|�������S��kd��<35�\���|K'����Z��LlQH��}�3�W�����������<�>2��=��vݹ㫈
�nF�L�����������H�h0���!n�z��qb��Zp*%	����96�Κ(��>��?aQԯ�Z��l$�u����(}&%u�PG��@��Ύ1�����
7$Ķ��(2n�E<H�17*����^@@�Wo�p�%E3�*�l����!0Q���@�G&N��}+<��P�2Y%g���J�~�Q��[W�����T<�;� ~,�
ǲЇ˴��[�{�X��k*%�̩�@�!��� ��g�/a	��2	��
U9ݞ����G�~X��3��L�| \su�b,s�O-!�n�[�A@q��3�E{jb�s@ZqF�;��@K��'��n��^���XofC8�¦��c���ҸA�v�l�I#���J��2/�gśoP�=킅)h{+�fq�oG.��NڪW�\��/�~��	h���mVH/��� A�O����TX:���U'���Ȩ��h ��mf��D����T�G~&ԯ�B{���6�����4}4� DYzF)-y�Z%'���s��VE��[�S��!�:��WH�.b��������M�)���%�|�`��M�i�N�M�@�'#f��yB�`���c�(�����5BI94��zf��&���80�K�Ec��E$w�ȟ2)�O��G�{��_�8RXTE��W�b����������P�����L����4o����[�#C��a-�������M'���\Ì���y���xj6��-���ܥ͢ĕ��ȑ�BU�2X�`�=%#�{X�!p��C�tnBl�H��� UId����,g��}$@��p�8���Pb�8`�(N�L�N���Fپ��e6�u}||�Y���m��߄���Ӌ� 	��v��$:��9B��x�c���H�?��Ps�&#*�����{�����?\Q�;5��2����;�lٶ����6YH����'�;1ؼ/��]C�7o$�@�m�X^��Vw����C����g4�rkX���ߝ%yT��DC�6 -������#L;��s8Z%��B�# uy��d��Ug���Q�Y�l�1��w@H�ڤ�C�oLdq0g���9�~n�Jh*�j�V.���I)cLu���m���A�kx6	= ʦ�X��z)VDQ0 
[�+S��09���ՕT�ЭxO7(���椖��?����l7���3�6!@F�=�s�p�S��p�����-Ç��mBex�XN
º��8"�8m=ʸ9 �NC�C�W6г2��C�������F���ba5+sA�L��+ ��c'�����g�=r�Ɠ��V�x82��̕�*��Iv+��n�˓���jT���o߉r��[�����s��`�q�X���,�%�ʷ-���P#iy�ƃ����8Z�>��I#�N^��;�p��>�Q.E���)���A娠�s����kճ��-b$�tHϝ'&2r �Cu%"��ؖa�k���cD[�P��A��ݧHI��EkѶR2ַ�&V��Y~[�U�Br��'аE���p:Q|kمM��Vf[r����Q r#����YG������X�8�I����S�D�?�R�&x�L���}IY�����3�w�� ��s�#
�?V�i�����x�OPCvǁ�V�Cɺ=_%���nH�Čx��q�E�J��ǈ�w7إ:ո�OXŬ�cV�W���QN��
va:�s6(�Q�?���O�q0O���D�Kr\im�=��!Dp��m@]���{��%��	l����bi@˶A�M_�kK���U�j�ؑ�u��+;���Ĺk2 � @�J�}t�y�+�­�����0|;����]�v���s��4X\S��I�i���P���[:����-���=	jϨ��wu�4F���8�0�~ѪD��炓�B|�9^��V���eWU~U�t���n%�uq����'��Q��`�{:�8)�.Gqް�������P���D��UYW�뮔�����6�^uIhE�/iP3<�9�/�p�W��� ��A�Lܓol�`	�!�$��K�[~�}�rЎr�9\����P%˼h�eY����i���CNQE��3/4b�I��`E���}8#�>q5I���@�s�?l���<o0��`���F���?Z=��3�u,�*o�<O��`���	h�f}��7�����uD��c���2Dg�s����Dx7[��
G�N-������k�[L�J>��Uho�,�"��g�;�M���l�6�KGU��&b���/�, �xЎ�9w��~�Y1[a�m#��c�� 	h�BC��d�W�:L$>7ڂ<�f]x��¦9���M�8~O�FMm$e��L�� ��\ϥ$Kd���s�
�	  f&OM7Rb��B�V�g�v$Qj���5��-/D!��W�K!��73���5������ q�@-�0V>;��P\J�75^yE��X���F`O���7�E��A֚c���8;c,��Nb+Ч�� ����V���m�]�R^6�U�'G���=�%^`3�C@�Ou�'�kܭT��67�T��_��b� �>Lm�^�[W+�[��Q����$�M6��L���C*�u~ԱXƅƖEӺ���i�V0��:@��(��b�Xa��vb��*����$��nbi���ǰ�+�����_w��*/�o7/T�་t$�W��C:��Sp-�N�.�fc���8�	��H�͍+2ul6���tj4�^ZP���fۼ����u�L����6�C��T�4��\B�
	'%6����Y�n��A7���&.�	�N�S�Ok�� �+Ʀ�9.�L5���l���"G*���F^��b|�\��ĕ�����6��^k��q̼c��i항�`OT}� >��MZz˳{H=�BL	���P�K:D:�ң��������!�b���T �sm�@�G�L�<<�C������,���<1#債j]rz��֮y�H@<�,�������J������k���#�EB��$`�#�[D�m�6O~�Y�$��2j������@�9N[�}����b�c�E�@Ncil���A`�����������R��&�1bgK&NԚ���ر$�.\�sǂ��_#�cM^����2�HY꼉96� \o1%q.�vR�+ �	�k4�?�&�x_�,my��I=�H1Y�;6��甾ͅ
��0�ƴ�0Q��!i2o���6]�f��n���2
/���������������Z�����~�X�':x�U��<unǤ�#0h(ꍰ"}m��.xޘp���c[I6'Z-�  �G��$2����x�R���zQ�@��F麻��w_�*�N&s��j�;��Q�w�כa�@O�����s�c���4ŤG1��JL�?Z�eg.�V��a��m���<)Pʲ56~�����r;���`�V����h]�ˡB!o4c�����ڟ���'ꥤR����.�_��~H�*J�o,6��<��p�c'�Ӵ�䆏q"��.;0�T��7�PqѰg�;8ī&�Z,�Ҧx[�j/��:=4�������a�a��m���&=��	�\к�:n)p�.�(
xE?5A�ϝ����б��Q����e�$A��""1�ΐ��Ϋk)y^�աbg�h L r���N�?H����}�D���վ�f͖u$&�����3�VL���	'�$�c�Lmrm�?��ӵ~��{@���xM\����X_k!�E"�;�5��Cyz�+���	������%i�q)B�Q�?�jB���o���Ƕ�8�Ԁ�C�m�tθ���k����@7f\�h��7�1F��v)
-d��W��Ug�1QFxb�ԁɉ�p���'7!�M��vBQK2�����#=z�a��m|��)�!��+L�]��>��>z����٥���@�<�_�b�euNc`�x2+{þ�\>��n�0����'P���pB/��<�LE8&��1MӳL�_$,�5-c/�O���W�ۏ��v��䗊�w�^O�J4(���l끫��2��@LD9۝2�]A ��s�͹x�U/���gU�C��60З�=j��LoX��6��1xb�U��^�d��G)�"iEg���iľЅ��)�b�4�_����y k��ς[�'s֟���Z����w��c�5�6˥�$���\��J�f@ꊉ�X�x&�
͡#Cl���H�w�s]�MbyzR���90��le���}�dt֠CqSޛ�i�|�'�ܝ[����x#�E��+��i\`��M��T+��n ��(�d�@eP?f���|�V]3���ԟ,x�)ܹd��T��|h�_������ѭ@��3�y?x�=s5o)M�.
���7�.�dM�]��9�d� t<큑s-v|�Wg��z��#��/.���?��q9�o�M	K�kP�t��C �xZ��9P�(V�O��Qtde,�O�캏���#j��ܧ|��:J��d�wf�gh�
L����!쮱�v��᫘�*���a��r�����3�W�U�����H��׬zH�P[`��鞚��*	t��(��3�fO�s�j�g2xO�L1�1|V52������C��>iʟ�S�p�?��p�Af|�D�c.��o)X,f��^
��-��#�JXŨRo<��7������'�-1�|��Ig����~�Q� e�Z�V�ǜ�A��pU��(9J}��Ø3^�5��
=�-�v��Dk�q���lj'0�X��@q����'4�����ٚ���2}K���G���,F�# ��n��[.E�e���e�eE)��]J�w-���9hx�Eu�>sw.��Х�0�X���;���%���bz/K������;�$h��ѽ:P��	�<�w ��я������t��E!�6������g�0��J�_W:VWP��O���+lˆ������'�%�Iy�F-ֈ���gf���U^���W�\�='�~�Js���	���,� ���M`��a������<Q���Y,��ETKu�K�rj9��,js�i�^^fJ �6���1��NT5�{˅�t�1���uλ9�cp�~��ro>�x�6��l��'���n=۵�_����/
@�'�؟���V��q&ywz���8�\)pt�"�>Q��*��	���+d<ƍ�|��������ľBѺp�-X�V�)�y�p@����[ƀd&n)���6ʱa���A�QOi�pӒ�2����1��Z���MJ��]̿�!xҤ����>�<���ˌ(�ц�xK/���-i�P��Ŧ\9�[���bӜ0!R�e�O�Y{�t]9u�t�v�+=\&���,�QW���8��L92H���~�r������ۇ�}� 8q�~��r�����!�'_�j�
�<0���=~
�ݔ[T^y�Qo����q�3�N��.�.�Ϊ8�WKI|UA��im@���a�z_�nzi���r����g���&�\l��=c�pG�c�%�	n���i�q��H�yꌧ�Jn���ls�uC�)���i�1O�O~C�JЌ��)=]��zF��<Tg�o��<#K>LJ7�o_�˕kPJw��h��<}W�u��"x�|�;	<��ߢ8gV:{�����Z*|f���ӷA�4��ۜi�x^���3��V�����'���	q�rb��h��f�$A2Q\��Hf�X�b+���u	�5ޔ�ж
+>�᱑�M
�~I�ͨR}�S��Ew�����˗z���%lDF6 M��Rw����$0�쬋g��?���4G@|0����/��vFMQ���%��oF��*T��R������zҟVBw���	�����I] �	1�iTT
R��A�/E����/|��F%K���w�F�i���!�.G��; &iS�x͒�n]:;�q��Q���a��)q�o�12�!O��ϒ�"��G���|Yy�T$����!3x�5{�bi{�^?�a�OS�l��HD��U������)D�1W��S���x+c3��~�5Qhx���ߖ��Hb0Q�D|�������.�PL�8l�FM�4#aB��q��~Z+V�bu�V� �������6Cv*�G��O\Dr�I��_@B�b�}��%�D�@�hC����re�:�ɾt�vE���]=�</=�$�b�כ�b�= ����=�,OS��F�-f�  BȔ�W���?{=�-�E4r��'��-j�亦fO�-� `L�Ou�gf����-m3%g���<y�K<�&��%��#���������HW#`�*��#�yE��YJ��I[��I����~!�{X��	 ��ޓ��z�G��:�x�R>����q|c~�#&��0+��O;qI�܊� �i�m�
���L*��#t�9-��A梮�3g�9;P���9:N�$�dք3?̔����a�a�4VQ���z��?z�c軠 5�ɡ1�"J>��a�V\����*z�j��N��Hz��r/?"�\�ߪw��.�9�Ey����Q�(�_Vľ���o�p*,�=���]h�2�$�� )�^��@[��)��z��
z�~� ���
n��`���#t=���Ow�aFd0#�~��.�h$�u ��ߨ�i�rT�G���9n��Ӷ��E��eg)z9q��������D���4��qZ��9(_|6���ȵ�0T;�J�j���c�|�&8GFs�|zt���z`F&�\2znoN��-���� �4���y��q����|
S�4�3�XCie7��8�M����.���ۭ?�ӓ��C��>ȦU�;������w�C�?j�|kZ��#DЋ
�6��
�S���9*��l+��� �Y����۞UMG�_Y��2ͦd^�����Զ ՙ�ؤ؝�)xo���TN��.+�O�Ĳ�h���CY�H\�!E�x/�������9$�U�j0�c��n��Od��g�,䧯p*8ȹ9�(}/J��������v��h����ia� L��|��4�u"'z��Jz
(]���P�ԝᐑ�ek�����ߩ������dv61�í��c�udI9�	��%h�~GG\L��w�$��y����ε�b�ű�����]�E�J��i��B+
ₚ�꾴�u]E�Eu+��q��!����7Y�G���A5������l~�^a������~ s�=J�5�d�Zk4pu�U�K$���'�D��ߕ�PO1@�v���h�u��㑳M6Em���yD$����N�̻s�?e
�ZZ
��[i�%��_hR�|��� �3�ەq/����(b�����Ʈ̯�	�7��)vC��`����� �jb�е@���؎�L�;:&l�.��J���sM��CX���������U�3-��6p�]�b��ݘ�v
 bi�:v+tk�7�
�/���2��~U��`>�1��#�Ǭ�!߳"�B���i��d<������ـի�o��������R��*�@�?f����6u��
J�&��v"�fjJ�e3Ick����0�[�5��w9����l	�T[�2�����kl~~'"�^ ԁ��{����!�e☨�	��o�J\���ϯ�6ꏚ^2ʦ�ّwf����S6�s�����U����,�����$��W���gyX篢'#��<�A�iT�X�..��D({�i���'!���=�9��Q���m��:�-Fb�A�B�F��Uu������13*��N¼߃(��wAؔ�Y��˶]���6:¨\bp#���``$L
�w�Z�i��>�k�f�(���͡���][*@<�{�<(�gp��b�ґ�-��x��U|}s-�h���! �,D�|u���ǹ�q�������c���M{�����>Q����4~l	D�E�"���y��D�����n}-j��tT���z���cH	��p8#{0��������U��oI��'y�%��*(
��}|�iʂ��]iWGX���g�u|�M�+\�e��m�L�$eGS��͠�� ���ر�;m�'dgS�7�8%?�* t����Ri�;ʹ��D.�k��N<�{���ɪ�{�O۰�@-�t"��&��Z);n{"�b#�F��e�^�FA?�2@���bj5��4�b�NLk�om�Dm^kޯk�E�^2؂y�9�7j>J���;�h�L�x1ά�j��A��DK"Y���i�V�6d���!����{���{8M�ѵ�,�,B�{���j����c�˅6-2��4������U���Nv�r#����}�W�Ac���)zW��Ĥw	��{�0��ܽQ�Ξ��Y��P�R����^j|oΦ��2��I���Uqf�p3���^^w�j���#*]�#�?9�8�������J4U�\J�;�/���N� Mg�[Dj�WD���v�Ak��^��u��m��E��%<0�ӫ�~�u罶��!tk��sa�Nm�����������1E�۾#W{O�_�`y�/��E�q�Ӂ��+(�f ��Jb�^��ú=�9NN���Bq��n�T��u��b��� �BJK����(��X�lo0M�u���sXXRr��x���]��gUš���pd�deL�����|f���@�۱9���c@��=Z��J�rdR�W[�N. �d��tQ� ����5�����8Տ�5iz�Z�=��q�֝�0��ٲry���� 9�?�S��[F<��Ɔ�^�~����Cp�/�c	�}�~3�}�ܯH��y��I�4��L>��� a����}`ńw<:��~vx#��� �ݠ� 2g1�&��T0��mF.���pQZ���1�v�AD�1S�[0DvZ_+�{� ;��a!�N���W'(��(%T��~_����9��ߑ g&���D۞�~�&&�]�)�u�/��Q�+R�n����(d-Dj��'�4� ݙ6���@s9�����/e�v�u���X@qO���?��H�3�~F�b6�eʨ�a$z�^���o���D�'��І ���ZE2�1��jWyGP�M�u&�ѪS9@f$p�Mma�{\^	wNşN#F��
eJ�� ����e�`<�+[�����H�M�9�b~�F+�X0����� }��T��3�}��k���h��#თm�Ga`Z� 
��LN�:��������������QO1�,5yʻ�Cir�C���ܤ�V� Ɠ����2����(4�ی��Ok9	�@�6V�2��M��������ȍ�膗_!d.� e��#Ĺ��o�*�ͺ�"�a��s=)9�j�*��*����m	�BR�����{���?�R�l&ư�C\�!e�yx�� ����@��<^j?��(��yQ��:�S8����"ɳ�|�"I39��_��hܖ9���9��>�_r��^�<q؉��~G��K�u���C�Zc˵iv"Al���wa���gg�	�A7�`��Q����7Cn��L��R)m<?7&��Blӳ]��3^p��Z���>�1!��с| �Y��e�]U���$��m�U��=���N�E��u�wrФ{��T�Ly�������q��k�ӕ��t� �=��"s�(d;~��]�i��2̠�-_�B�chE� q�'��4�3|�u�@�Z�re6�O!o�#	�w����_LJX��<����Jn^�<��i��\ߧkB3�E+<YE���'��H��>�:���3碘��n���x����؏�`�8=��np&�=D� s�>��^\�U���1��Q0Ϛh9�y�Fw���/%���i�1t#�T�Gj���chbwO�T1�zԢ�L�4�����8�W{S��a'*ʳ\H2+ze��S'���H},��	�Lo�}��V���~��B"w�+��|j�PeH:{QJY�RU�l�nȦ�?�H�Y���H��k�`z=��1X4�����0�!�b��Q�I���nc�'��æ�_QV��v��������j�����zW:�N�h�t�	�R�"F��/�$����u�S��[�(���*u��]m��� e��"���� ���V8�N�_H�	p��>Ӡ:�d�0&WElM���n�_*&�$y:��=�X����Ǉ]f��pl���ή������� T��*��e@tI�Q�2E@V��6 Z�_j�f E.�aM,S>���E��4d���|��R�3��N����֊�MX��ۢj��m�1�\�]�m���qg����`�� ]ur�Rأ�A���y ��SG��DC���~KA}��PO����y�>���\�mV�E�����$�W#�s�UK�!{H���I��#,Q��#��B�2��	:� 
�?@*�X�r�\=JFz�=2���6\M5TJ�e���PC���g�-k^8NS_�hY�%c$CV9Ubh�-0k���Ľ��3�GR��� �J4n��*���@��TqZ&�`KK&)�������}H��-�c��Wcr���i��ւ�,�~ܽ7�X�..q6�}��_aᐻ��?��1�0"��u�ь�2&q��߫!Rl��"Fպ���y��y4�����#�(��7���"�<5x��j�R|�3�.�Z���'�[/
k��t{2��+X)��\d�(�:"yS�	H�Q��G��ɢ��h�<���
&?#[҃����3;ε��G�=hfĤ-A�G6p�j�u�I�"_Τ��A�!�a5�'T@ ;w����eT�:
���|�K·��Y+g�O��i�?|ypt��r�?y�U�}>(�;�W��h���w� ��M�睢A�VʕZ�n�R�r*�����%�D�eK
hU�� ����E�Ț��?��|�Q�j��pz��缾�L�E�Ê�t<���Кw�i5p#G�&
|�a5��Q�j�2�m�.��U�]�Q����Ixs�H"Y�%f+.�"��)^�bƲ{���.���i�%���=RA���@��xv����B�1�fȃA�����;�H�ż������AH�i�ogps?�����z�z��f�l� �Nvuv��(��wIl�ۥo�6	\�'̪���S�5�bK�H&{8~�"q�1CF�z(��*�+ >�X�	��D巆؃<9<x���^!':�fz~d�5�d�ɺ��N�l���0�����/VD�u�kϡ��~�?��3����#l�>^�9����r�߭/�Z���ם1o
�����c���0�[kp��x.#�r�ɜ�j�����=�ëA�\1���BRY�)ڽ��	}��"��U�u�κ��#�s�j����p������h5R�c�:Q�:�:6�yV�S��d�s&�!7�M�@_fGw@�-�%2����a9�=�3��ӱ̔Ɏ�u��B$+b1䑞^К�H��O{�+����"��@�ƲF�J�	ލ�.1w[����^QJ�*6�!�R�Ǚ7�좐�: ��e[x�d�9�}��q��05�Z;�&�2��pK>�{r��>N������*�j(W�N`E�7& K$�1��r���C�����a0�A�fe�bA���+@��q�1C�����O�1�<@x��6��$;��Q���I���wkd�B�H�؈�LYi�O��ɳ`��&�)8�|�qK�֨Z%hǧ�Τ��}�iJL����@6u���"O�����.+��=Qayt,��T�ˍ*�\��i�S��f���z�Q��^�m�YCxQ����Zo־��$�CsI�C͠��*J����*����(Y��\<���o :!o[��eGd��j��M�� b����d�CP��^W ���~�a&�*�02��S|1&��۞��T���A]���=n2g,~���������Ĭ�#^1ڈ7f�a>[���[���o�B���� ���M֝�,b/���l�pt�Fa���O�"�D3j�#�a�Ĭ�����usf��$J�/H����e��1l@UE��`�y�r���b 1��
ɤ���,�����{`e��݊S�"�l��i��N� ��r��ψ1ap��N��fݰ`I#j��+S)q�SNǫ�r�8�al��c��4��w hdI�.%�?���('u�Ns֛��9A�d����ֻ�|���xV�B@&�I����LF�vS�#�c�F�n��|!�F�!����1��5x�
��gv唣�軦\��w+�BG��=�2��J\|����^Ŭ��^ä�|�x�S۝�%qH�c}�0�t���t�\��Κ��ߚ&���&#�;�2��+��8Ͳyh��LZ\fˑ����g7`:�I`Q��nyE��7��-�����i��e�,<���(�PyL�@z	rK�W���Bm���4�6e���gT�:P�8qG�6�D��T ����8 R�N'��D&�4[ځW�.iF��F���5�B��k��~���,� xd�W�BS��(��z��MҾ��i�꙱����/P���}ӱ��&�����Js�:3xbIo�Y"8 �0I�&T��%�OS��#f?�'^ms�����c�L�>�"a �Q�Y�t>�u��f��޽%��E䶃=s>�F#3e�B7w�ʔ��qN���9L��4y|_K���	�E�cƕ��������:uؓK����C��k�ԗ|x8��F�%}-����2��t��H*�*'�QԼC��
q0}�.�<)��� #k���Y�|��V9��M�\9�H4�����o�AB4@��bk>lJ-�����/zZ ]��<c7���:�^�;�}?�0��V�|̸�+^�Is��|$f]7ʫ�R"��=BG���"�^�>�g|V�ͬNL[��G1tu�Y�s
y�M��n~2F�_*O9�*!9���c�y����a֌[j��2(��2�(��v6e����k{�N�#�>��`z���`_�,H�Pk�%�ul�Sܒ� ��)�v��g��;�_�0��c�Q7ظpv\LN)�U΀V���FգΡ�j�)�
=O�������f�GjF�\����Q�g�vf�C�X'��7B�!�n(��lo{ī�L/!�v��|�,瑴�\���[�')_[}U�8�B'��E�bbdyZ��@�63�T-^���_�׍�?��[��C��GMA~e��tEK��\���b�@��aaʱ�P��85�HAщ9�.b��a`ʛ;�8m'g'� t!7&�g;`�˩>(�'���]����.�ja&�䢚E�j'�*T�j��[���+��XWa`�6PE�r�@�U��a�+=H�A�Qc*������NV'�}&�$��]�!فj�|��hB�hs��f�|���|g���-!�}��
�:W�q�.!���N
�>��@=H�H-yig��Lї%U��=��YW��	J����{S��u?OE�S�UDSPRB���w#u������U�����8G��E�TOS�����Y_(2��ϋ������|8���YڂO4���Z�N+#	��Jo�Z��V)Zҭ�} B+��N�R�
z�(1��&���k����ʦ<�=�)�"�c�I�f*]I;Є\B�'B��� �(� ,?F+I�S�}��4v[��K��Ј�L�a�M��
C�!ߣ�ҡ��"��w"%���n��٦'m��J ,\ur,-Ȯq����Dъ�t���:�Ѓ��ű����|Ґ��믓�I�Q~����'y���+k;������
��v-ӡd�?C/.A��<�9o�`�)�#�1|��uJ�m��ّ�/�h�8υ���Lߡv/b0l�K[պЋ4��4�l�^�f�T�t�V��^�-���rN���&ԅ;$�6ձ$*�f"K�u��B���K^i��s����?��o
���r�]��h�y��[^׾��~<�S��t�hɄ\��h�`X�x>�n��)�g!�`�J.��:&Ѷ�]"0��!wm�N����K�AC�	C2'�x����k������&������l��&"�#�b�?��kB���,;����
]1��i�SY��\�񬬩W�"�b3�|�`U��\�$�a�A.��/x_�`��];7p�Jn�&��(������z�?�9ӡ�AU*��=i�a:������$�po���9�)�0gOC
��Q����͛μ���*�VӃ��.��ϊ�k	ޞ$9�z�?U���<Q>�dn�=��[�q��l�'S����5=�q|�9h�����Gl��#ѕw��dH����P
�?!�s�1���y`n	��~��®LK�#�GEV���r�i^�q��T�<�7��ܵ�j��y�cX�E$z�����8���E	�!�2�����rux�r�i�>�������}��+����0�,��8����N�gxPd�y4��ܔ�)�a)_���(���G�� ���R8b/�)�A����Χ�z]j��n+mcwI�����b�ś��f���=��\F�I��18dh��7���6�4Q�x�ek̭�5�[Oӧ{�u�D���6�k�.)ZW��
 7�}���؝H�v~.����$�ɫ�V�E�#�4kJ�h�L���W!� ��`�����`�&߁�v��0-�5W��AS�Z�?t���i����<��"��Ͻ�΃�v:�S<�����H��0����7a�<�"O9��1�3��{G�(�	-)�p��r��2G��"��˳V^����n�3���q��K������Q+���n���[��j�`�E��Nf�����d� >��]ႚ��0X����U��>'=oDp�����Z9Є�j	��Y%��|Z!�$ބ�����{*^%Ba,N&�c�Df��ʯ�k�u:=LAS�+����&û�4�/4:�L/%��a� ���Y�À��u5L�k$�/��u�ɷ�D�!�Z��i��V�W���bX��O�u��:ǧ~����J�ȹ���ʅϥ�A����$�FċT�K��"u<|���X�Ë�������]<�� ˍe��=eW)�b�EG����o���RFg 
@�~�s�azx\(�5����0%q֣@�P@G��b�kn�1��T���
��{���E:_��V��k�L���bb/m��0
�;ǋ��WvM��;�_}Q^8G�7����Ws�͋�E@��L-�<�zi%����fa��k�D�vL��^w�>���yKH�aSy#�R��Lqw�	Z�}+�cÅ��c �kD��JW�eܜ9U�x�$"����Ӳ�] x3���p,���I��T�B]�D*�%SM��u���vpW�����8����S-,���ؠ?[F���b�L*��뢬�r��;�&��^��,�yo��\O�`_������N�V ����,�6���;h�x@�ݸ����j��`�yq'�ZlW;���M�/��(7�!��!)����)�����Ae�n�gt��v�����J;^��ج�����1�0_U?�tᎃҟG�A�L�52+�xS@�R�������iP�Ϊ���ȕ^�ڧ�t;�{:�bq�fY�ō��OA.� ��z���#/�ss�]Q�nH��2m�k� ����7ރ��$�y��#)����r�������\��$Jf�"�M�L�-��o��9�Xh�X`=�5�yE��QZ�Sʹ� F�_��x�Wc-#RL�3i[�(�����=�ym�)�<:Z���|I/}���Au�g�8xk)��		d`��y�/���[�=��\�q��5y��V�LS�FSA~m//-a���c�{����ϩ�c��E`����#xoi���RL;+a��C
�L���mea�p5	ӓ���x
˃�"��k�����Y���}ab���BQ4����|?(y1_�������nmj�^���&s�(*#�g��0������ա`��ٙA<�7�ۯ~(�7KZ�Av�
̽����o�{�:�7�p�"��si~�@|����d���'�pL�{B L�F�B�RLrƟnkű;�
�ɓ����.8yn��_�i!��z����Ck�F�ʾFQ��'I5�� @���I��a��,ݵ,y�oݙϨ�lwaH�OA�����G%���Q�)�4��Q����s[��`
�������Xz�(�\���aq��c������%��['���d�RR|�䚭���
�u�H�$*E�$@�J����4���_5~��S�����|f���� �#��Sgd}�)��K��;z�3a4�݊�O՟�T�vƅ#�&��<�/�,����I����.�i�?�6�6VЪ�=��x����
u��e���{���Xw.߅њ�����0i e�9!�k��|�6�Ỿ̶��{Fxd1��Ћ��Z@����5UN�<I���Τ���<����TÈ������Polo�%{{�Ox���a2�^Sq�i�#a�?�L){�{>��h���Jg��l�"Fԋ5=�
j!�W���=��@mHbw3���M�ŵ�稔����~(P��'�}���a�����}'�6��M�+��O�z[��Ƚ��=���fk?B�cv�<����v��=�*���Qn0�xK07�͡d?���l�iJ%�ʜ�z��|�!��5��7�͉=0]y�! B�\F�;��Z|�N����Z��Oo}�������?4���E�#@�`���+R��e[��-��)EE�Np�{N���f�>�l�RfR��C�5n��ϨK#�����3w��ر�z"b�j��敊�etwDM���t�M/�C�6gD�����7��[��:f0]�V�cn�V^�!��Uuw޳bA';p�E�ݲ�P>���D��А��3,�9a�q�-����"���蟷���,�|�����Z�(�G�ϻ�����(`���n���m�E��X��>�4`��UȲ���q�Pܽ�
��O�o$�� �Ya�D4Rj�<�}jڤM6|y|�(ǥ��1��?��a��Qbv_|Kzk�47/��jA�gܦ��")�L��آ5J�%�0��U��̙o��k����5��Nj�;p����h�ݮ	P#~|���2r��ϡ3�6� rD�"$O�"^����?c�qo_��K�׈�u��A������7�����=G��ߤ�l^�U�9&@���0�~��M@>�>8B�;�%�1$ބ��M���WP�L[z�	u����D�З9�6�ɤ�>�ʯEt(����F��q�p�;����3�#�s$����z�5��OhC0C�xWEK����E)������1����Cc����}��;zK�JQz��/г!�0^SBm���p�>�H����1��*��p4V�E���^~�V,�ʢR*@u�a�F��	`��m�ǔ�+
<%�C���r�����F����BLP��"|�I��� :nZ�T��u4,�NΡ>dוՎ����i���"  ��3�#N���M����Q��Q�su�:�H�.��_�R{!��u�n��D��{,5p�r]avM䯏5%�V�ɞ��֍W�.e^�d�C�����veq%J�ӧ��&�S�*Pjq
���Y�3�Bq�Q�f(��Be���E��l
m���
1�}z�r��>F���xqW�;a�@/��`�ь ��_	������$}ů���|^�NiC1ӹjE����N(�8h�M;�?���/>�g)��=`�u�%�1���_Fdbl�1���BDW�<��|���d�=�I����G+�f�zG���D�l��^�e�~�|T��ƖƲ�^}����3�}ʼ%���1:�PQm|-.�"}��H��P�K]}b���.�Z���Qo��&�ۀ�f-���2)Z�jz )h��B�J��tB ��-�>�M6�|��$a �q����O=�-�"��O����>Q�� (�NU4�{9�vA0���ar@j_�*WX���������<Y�{
d��{"--�΄�z�ke�������[�%�rOW�L6��A�h�S��B�%�5�j�-���/I{Ѷl?!tDf�,N��7@�a�й�kGNJG�sGYa�Ш	N�� 6+��:�$�:�Ӌ�����^�A����l���W:Ehi>HZ���>ba̼0�v���.��B�i鄂���σ�Aw�3�|�w�^Y�4��1�Ct�j�����4K�ã'V2����q�l������?@�ꛬ����R�Vq_�s�	�,�N�L�1[���'C��e��{ ��<�K����kk��W0���J���ظ�3�p��MP���]�W �NC��2�z����fm�>cE9}.a�3�9���{RS<���sC$��ad�=�>���\5��R>r��{�����_��*@�b�ZZH#Sr������^X��4Wq|��ѻ�P�k��BW��ԡ�ZNr����(���꒺� Z�+|^4p0���.�)��v�e;f�5�xK�����v�<�.���l�˻	 ��8wxڅ\2O�v�6G�Z����ZW'�h�����R˭�tXlͳ���+3�� L�_��cl��̾Y��=P���<"�����{==�aЙZW0S�7�젓q(��Rx�!���i�1�5jBr} �I��;Űy��h�Z
��!�ёDm�����xW.=�;!�a�;�������UE̓jr6����ɡ �󞽥��\�\�2�kɢ+<�FSL�п��7��d�|���`���\Sb���l����T/\���*KaE�+�=���@���G�	{K�e�:�Ga�{&�+X�8�-�C�ClPt=������yJj�*��{�.���s��_K��  ��fhq�(z��BB�W�~/�ϐ�f�BQp��~D���s�w��':!#�8Q�SF7j$�iX�A�d0|0�TZ�f�ɬ, �G�q	?H=ư7ak�q��H�ɇG�+.\���)�/�F#���S��y*
L1���S��o>��!LOw�%l��!��.?�+��Y*����1��{�}�μ��"�k�ד�u+�-�����dI�ln���wHk;�)y��y ��O"��PJ�$��_eױ@�#�0���P�J�O��P�]�& �48�d��fa�E���Y�җn��U�G��۱��D3�s��qϫ�34c�=��C~7�:|@~��ko��]&-��B�!��%<H�H�`aߢ1�U���I#n��]&0%�n����9��Ery��2DʨM%pH�g;��b���Ie�]�.�l��v��}��AO�f{�6b>ݒ���d��^�Nf'�L W�F�a�uܤ���`٣nG�׍�qd�E�2\x���w�ۻ����&aTɷ�fSѸ��b�T�+%6�~��9^
�s*s�;��)����s��=P~�:d�<!أ2'cކ��5^�4��������M}��3o��X��L����<T�Aϣ�80��^���-Ρc�X��������N�xF���_��ׄ0���B��7���;8�- >J#��?)��A}*�����2����&V�um��w�)V!�WX3P�rb��tl��rn`���r.�e�g�~8ŜoO59dT-��#��@ТE��p~�`)+�}�p-ɕ")����,YF�8&�92'6|�#���Q��)�ђU|�0�p�Y��B�*��1��xq^z�#
`*q]��#�@�fv	�%� 2�u����PY���b��`ڒ.T?�?vXàryf��B�fm`�y����<��F���� ���JZկ{�K�e���I9h�g�N����T# �[��
�.��t���NL 3>���C��7ɢ2�j�������~��Q *�%s��{(@Ƿ��2��'	�d&W�=���w�d�䉏�����$�Q�)��'���s��D�WL��7ҲT:��!e~����s��*� �Oʑ|��������Z�[?����I+�n��7��f������4l-8Hd����� �5�̹l���2��	�E��>M��2g�I`h2�e<��W�!�a���u�JIk��mxϙ�>�K���HO�iR��#��������̴QVơLѿ�Sb�N���P�t �"��HG�F!<��(��bxx	0 ��D�Z���Η$ԙw(����a�TI���$gؑ}?��ied�\i$������6�/㦓�;/������GƋ�Y$\�{�Sl�z`�.T��ז����o��)@� �N��#���~���z��ƞ�!f�Ĥ5����{����U��;�/�/G�i/܄�G�c
�{�K�^�������a;��l*����t��2_N������AX4���d�P�6����3�]�Y:��5+Z�$	�t��.��6x�P��F�f��/ڛ=q���O	��dF���xW>����gЭO<~F���d:Ow�2Y��{��JaF��|Mz0]����ՙڕ��姯��B��Y���Vn��_�zD�l!ʖFs��[Z� �	��pF�gTT1�nm��L��h�u-�TUAy�V��D	^Q����A���F����<C6��fe$.a�o`Ʊ��M�I���aAu����z�?�{��({4��߻n���lH��ٲ�w�V�:jx�A���Օ�.�.xc�C8L�g���C�M�`((���1�v�����O��6���9E3$�{��z�td�{a�q0+��Փ�0�?`9x�˄��zv���q��j�QbLP�ĄӬJ���9�c}%��P�������� -�B�[5�R���g��z�n���[D���$�YV����R ��Ă�A���u�r#���N��aW���eI��e�P,_�꒞>6�ƹL�b��h�aZ�E��e�U5��=��1v������r�~���M�A��\/�	&l��'��!�ˤ-�=x����a�'-�6C�B�۫V�������9ZD���J�`�줒aFj)����+����/V�Wс��Ś����|��g�>D�Q�w��?�ۼH����Y���f*�ۏ��2�w̰�i�(52���fMڴ�d;2�y�"�Pz�nΈrœ\���!^i��Ψ��~�=T%8�ę�M��ʈ0nR#�.��lpP��,�F��0��.<�\jM���oci'�>��*�F��|�{�}�e��^�c��a�g/Ӊ���A�B����b�a.ɭ�,h΋6����ɅRҘ糳p�@{��3���U�L�5E�����B��zqr�XS��M�^X��8��6"	!�E�cqV/�ZI�/-X�4�Q�t�y�~���.r���4ب�N���|��M�f���ӊ$��KO���Y<
W��Td��x�$U���xb��s�U�cW���>�p�Ձ.���E�SB�D�u���rw�0�Ug�(bڄ����`WoCEF�:�?O�[ dѪ��{���D���Z�V����$�8�`�3�9e�P�h���P��{i���N�xDk�&�eA�R�
.��V�2����ݵl�_�O���_NY���㠹0����m��ܱ^r�����o/��H6���#�=����?�	���xBO�$K��%U(Oߎ^����9�E�_��ٓ<M���V�½	b�ąkp_`f�2�Uf�B�G��������!̡H������6��Y��UE��RBm��A�6��W����z!���M
?�4�q�.*(�ݼ%H�U��e��ԥ(�BM���j&J2/�?���fg��沼Q=��t���X+P��a�ȏU�h��=�A�
�U��⸑N�Ws;)rO��V�����ׁ���/
�)	Uص��G*�b�"�"\ǹ7 ���^`w�ln����y�1]@�&�&)h{�>��-��F2JAGKB/�;��ۢ���C��w� ���S���SI$�A������{b@����w��b4VU�D�I����J��;7�i�� ���>�w����Z�p�. kn��Pʠ-�a�&��V�1DѮIJ12�r����Xr'������C��������nVp�^ԩk���an�!��NF8
�
rPVN\�?J�)��0͵��o"��s��Yڠ�{��?r2}l�@)n�.���'~�\+�T�dg9h��Bo�1d���.3T0g��9g���Ɵ��d$'��I�F��[���[�L0Y�2Z��7��'��M`���-�6�w���c�L�1�W���-�A�P�M"O^q��b0E��!�;��m�vr5j�xLA���������~nG�ե^0K#n"5���KԗэWi]\d����f��i��e:/�g��+��epX=#�i�5
a���Q�����'�竪���?�B�
��R�6�R�O<֗q�^�hw�[���V6��X���A�!�F���oY}���mS��\�jq�' ż&���\���[��ڻ+|c��?�\B��^�+�I^9������\�܃��i�OU�=x�w��X͖�*{<cֲ�,��tO!���B늁�YQ�ZĴ��?����y^3�H�ވ�~��/��[�Ar�f�X�������V�s��b�\P1��^vxmI����W��s��.yP�Stq�aO&�2HZb{�p]���	�.��� ��2M�-@#���!p�q���8�s���]?i��������8s�C�I&����	�����a1
.����@G��K����	s���nq���������#i�֎�B�1@Ȥ���0�{-��cC��|F��������R�|�*����u6$'=b��(���4^KOC��%���Z�e�E�[ږ�M�����&m>�|���X{W����j��J���Qq� ��m����
?X��Lҫ|Y��a��y��A;����R?C��B>� .�#g��V U�V�}uf�B�$���YH[�!��x]3/ �d �m{��QX"::y�>�
E��`8�E�L��MXs��K����F�S�v��C���I���i��]�`�yԲ!��&"t��y�DN'D!���Չ �U��[�Up��N\6e"b��.�x�ـ�v<���XWo F��)>�K�L)z$���-cu
ox-	��*/-�YmC3�:ݮ`��l)-����<,)Ƭ8�GEBc��kd���k��ˬ�a �Gw�D)�f�p��H����a���-[hr�[-��7	nu7���5�N�w��ܔ�7\(u�O��h��P�1;e�7���O��G���&A<��Zu�kZ�$׃�Mu.��C5�j��-��ڽL_4jH9�Q��C��ݫ���0f�&FY�?=�\���0d����Bt�E֏����Ak�!��������T�7EfԱ�R�� #���j��)��ɔت����u]iwW��>b���7.զ'�cgI ��a-��(���E��Α��q���,Oi��̯ں�[���VMS4x����Z��A�PF��D�[^8;�'Blz,#��K�o�����N-�C��E������e��vHƽb�)v|����=鏛�NJ�|�W�Xt~X�w,��$�|���o�s��<��hO�.@����]Dvq궭!C�gp�x���>���kM_���	;��<�����k�2*�-�I��<W�D�Ӗ�/������̨*�/�q��tff�Hղ@JB����!�'Y�����ꡛ:xէ�[�����>G���ܡ��W$线��A��?O��2JL��!|,[�l�;!=��`J⋫3-t2��c
��m<�t��v;"k��psK�З~@!R��������x>b�}�K��#��E�N��J1^H� �E}��\Q8z6�a^�o�)3���W@׷��櫧� �4�h2��á<��>����&2q�<:�����b�i��F����Xi�W<�B	#�A�0~.�
pbg�	N�y��𽦾v�<�lW�<U���ym�B⨼���ʹ
�>�����
���O�٥M�З�Y;خ� g�\f=��KO� /Ԕ�q̼�Xb���(�4{㠥�oR�j>l���d�!�s��.#�ǬZ��4����<5	�%�����ng2$�����v�@�Ң(��]�F�Sf<%%Z>�dP����ɥ�Sç����U����~��&bR�8�����$�ձ��,?u�#a��U��?�~,���tŸ5����osB�5���[� ���#jp�v����$E��h̑C����%qp�m�|}z��0���˲L=sI�zL:��A�!����u�E�^@Wd��ߟ�������7?�>�(�L�����z�Mx�I�Q�aK3���5=���ة%�6�/Յ����ߞ�#�{��]������ow+g�0��:��(T�SЅ_�JFA���mNj"� ɥ<�y�'`���[Io��{�~?�.�V]m/1�kb���G��Et�K�^Z���a�y�W�U =���8?`���+��˷�]�<�C��R݃�������b�A������*�XftKw��%��ś�?��S�&f������H�Ps�(�j��s� ��K�h����g��v���Pa
)�8ȫ�{���+��1[R�'��?�[�%�B���B��a6+&���y�<a?���x��(����I"D��C�|�NgwU6(W�3��v���54�(	�Q�?��,P��K��<�����[K_c,���{l�_��xD�����յ���7����;9��.<#�����J��s1�ULN6{�Sm�eɲ�.�ʠa���u|p�'�5#�N�g��c������I:�7��)���?[�BFC������M�J�9~:�u�����uL�1��'[����o��[��hak�3�C�(KW:�V�.)R���M{EOi�87n&�0;#u���j�Uѡ!Qi��.���rɘ�����P��*7��\q��V(
u~w	U(�[Fq���^��ؙ9�Rf��O��Q��3j�*,eEW��<��k����v.�ڟؽ]�Q�"�<�<e�a�/K
_n�F�ww@�C�.��} %�	IAaS��{�[��o��$TE,+ߋ����6_�8)M �J�E!;��g����.,|�O1j^�f�Ⱥ�L�u(Ѵ�6�L����lU�������TU[4nX���$L�'���[3ЫJ�p~^�@vN��W�\	�������o)�#�`É1����\՝�-���R6r��R�Q�Ҫ-�����G�H�f����G���kVd���CY66Q��b,����6�/�>L.�H���7�	p��ZI��o�O � �i��켩��=��{.������/hyYz�H]8�9����¿s��~ѽ8��tQe��&����ؕ$Fx_(�G���M��H�+�6�P�/�$��q����X�ɺ]�S1�oPC�a�f~Er�x)�"�o�l�!	�=c!A<��v��a^��]i2�Fw��^:�#�D՟��H<&� �+(B���O���c�;]��8ȼ�J�z�u&��l�oL�d�2Е����V�DX�5#л{��L]0���h�l���\��KZ���w��A�������M��Z�
n�������oE=�!�mh�SW&H�ѩ�b_(�΃o�&@��/c�[_O�4���{��>~�8��M����`&���d�����y8��2��a^�(����8 S�o��Ήn}H� ?��^��
�]W��l(��$>#@L~k`~���{�)H�J�4�+ry;�a1`����i���+��lvI8\�?č�@@���~K`��Ɋ'O�{~�&9U�k��P"�c�Ee��<V�3�j����x4]\vi~���n���R��S^���p���I|�#�W�M�f���_�(��V@�N��Q����i9���:�9Sz��S�+��:e`��\F:��KFN�U��	ɒ1�.�_�Ԯ�s� ��R]�e�Y�߳�c�,z��g�Tr�>t��E�vj_��\⠕G�s��a]ʒ���t�ob[��ܝ	�o�?L_���4n�f���xȑ#;Џ5^\���d��7dEi���o��yj�i�r�0�G�p`���u 6k�P�el{6o}w���
%���0�E�8^�\e�(���\4��ژ���T(0���)�����\%O%t�5���P����n�k���c��0��V!v�*���0��w��W6R�a�&��!m��W'��Ջ�
����_Fo\z����</��۝#L�S�����GW�m	e6�5��:�E;dj�L�R9��d�2�r�7����3�lV/-�ٳ�BH�Px[6�EaU=I ��o���6�0*:|yρt�G1lV~�!6gR|C�eN� �/"�t����}%M�D�J���dSΛ��!a'/�J�TfL�.*+���d�2��m>(׫�=��܇��E���Hy��cڬ�ԩ{�(��xE�I���'� ;���e����+�@��N5�q�����ki�X�	��� �u���a�t�p�zɸe��O8�uƥ�=�Ӡ�% �[�!2�.��n�$>��J��/����׏���ϼ*r8���Ζ®����9&�xE}�Se�au�'�΍�c�4���G�˵7qT���i�,~`l�;����-4\\��,�g�v�E
>]͞��ɔʺ�V
��֙�ǩ��h��b넷Z	�<@�%Z���^��N�J%��n(���S�ྞ�Q��sa�G8��L�rt*���,]oڃ�euMĵ�o�;���	�2`��������tO�o�-����/�0Z�l;���%�F��D�vD�-�6Ō�vw$Qb����6�{�N��h$�G0Lr�7ߝ�Z	�{]	��i��7�h�������W�+�l�YN�F)@���\ ��9kB��Q��;*�l��1�}NT��3�v
�gqf��zzj��(�}��>�r2����i���LDA��_��Eq�c��C!	��,��W�����f��!�����7wt?�3���@�^�|wS-Ei7=��oPd�ӫ��B��ػ�G���/ �%Аy���n�;B~=���٦��.������g�)P�,[��ur�ɾ�r�������a�L���>�9�H`�<�a7���=|�D����1w<"�%Luڦa�j�Wa�\k���v�<�r��UU}f�Z	�"~:�L�EF��EI(����ы}
c���߆9RB�=�@�s�<�������<
�X���$��������F'���>m��޺_��E�Ys���L�6�=��CS1(���}B�F��)�J#����Y�XNz�53�7��oϛ�#������s��ˋ��䴘����b V3��4"h5�D�|MI^A��� W��p�Y�?��o���Qj��g��Z��dg����<��2�7������3����@@J��/@����g t8�U0���4���1������6�
9��m����0.;�\�RJ�{z�@��ƣ�����]��eW$�L��i�������#GnUu���������-�nM�Z2\^�9�Kй۬�\�2��.���+7c�����5s��mfB7?���Q� �;��������������By�U37;�j�y�rH���r�%��I$@u���;�j�9���J��׾�D[������J4��=^v�vZ�J@��N/��-qQ8WK��b�� �4���;B�iF+R[*�<���P��+�\�K��� �#�)E�Q]�<�XW�-T��X��y��@���elk5sb�u�E(W��ع�
�P8&a�=IOé5o���8A�T��j��_Ց�4],��4&x�*4��[�~�̵R����O���ަ��<h�0���!9ӴNL.D��x���m��<���3)|Ib5�UT�:[���ߖР�cM��.��.1����i���?_F���X�[���Ʊ��X��%J�������E�&~�O�f�2���q��C��
�����I���DH���7Gs��?2�G,���E*xSg�	�q���k�0\KN��I�v񻶋�r&=gc�����{����6��݆u[O7�ཪ> j����r��!J��l?��������q�6IŮv�9�%L.'f�byCB��XHWl&�;��Q{,ݨ]>�H�@�Ʋ�R���=�u���t��[Y�~i^����؍������G@5�.��U:�EŴ���֪X�qm""�EP_J7a����v��;%"̀�p�����d��6�H6q�R��n�4��ϯ~+�`�*�ID��dƍ���=�G�բ�M�9�|�$|�Ƽ#�I&3�KlVv?��UT,Ѷ,]�f"���b�c��Q�*��N�E(�n��j�ms��U��{�f+{)��q��S8�3{JӒ��E�������@�2x�®4/�wG����Mw�i;�Ō��r�p[cF�#�b8��[���LO��:�Rt L���gB>ë�<|���eX���E��|7��������^e2Y�Ń�}�~-�ր_���Ji"�.u[�[G��e�N �)ڥ���&��N+����~�:Yيq̨u;�H�S��K+��Nu���$r}�4K������� W��f:�<�F"2���=�<Y`�J��-.z@;$��f���{D%����3��h��_�6��:���"(d��=��_Ar��aE�����2�$G�&AP�`"te���9�{1��62��yQA��!�\&Z;�J�}V$�,q��]5����b�OGEq&}j�!!ò�B�G4�;cç�Hvk����79W=F�О_q��a����� ��'t���&�j��X�e�q-�1;5J}@��6Nx����TLi�ץw�C R���ԝys� ��}�r�����O�}��\ G v0vwcg���c�2в�U8�ntI�Q���8d�Ǿ�rD6j���~�{����H�������Ӡ��(�R�ٜ;潟�j �Re�7H9}������t�gC��7�Z�hÏ�nh��<����Vc�㪦TD�xE�APi����J���S�A�h�ZP���6��ؔ���3��_ey�A>�c�$��Rv�j���O��(t�n*�I9�؂h�-�9'�H��I��b6=�n��<ٻ�+���X`�8`�+`_�����镺�J��I�a��8�������>ӿĽn�T�$���CiLG)E�b@�n_͏w��R)��t�Sϙ�>n���Лz�f��.;ŐK;d*U�����{���β�@$BS�M��"L�1ݵ���1�Qe����Y��p�,/+:!��ݦ����7�'�K��m6����䆬y�F�M��$oy���x�3_���X^F6�O�4Ҽ��.(�������"��d��s�`��X5��m������Vm�)�Os�ԫYT�ȓ(O�(��~����o��+~�E�#�3�a2)ϐxVh�w֮���z(T���qe����mF�Nu֠إ$��. ԇ��Ʌ�S��g�����A}6��3�-�#�>��i5�Q
���ȉ�<ՙ�k�_ٓ�c��q�g�m���	�8��@�w���U��$Ѷd���q�;f�컫�[h��l�(����h���.i��(U�fy\%���S��Ĩ�s��w�6�$��ky)��74{�'V'��Jƛ��03 ��u����MBOG��׈ƽ�_�P2��&>�	sZ���ML���t�f�E��޺�_�/9f�w�x������^��%ؐ�"��#���� �vg���Wr�,�&(f��Ϛy��z�b��m�5�@�|��y`�e�jej�Ӫ[�AeC��ݓS����D(�Nj��(J_uМOPG�g#%��zz�h�s�	����(�2�{��䵧R>)�4����N���Rx�H@�g��d�Al�'�v��6��㏄8�i��`�1`�;�|�:	v��T�
>r5�BX&����ob���G�˒^�Z0DR>L�fxH�E~&�C$Ӏ����^o�.!�v����,^bm�<M�ψ��5ؿ���˺t�,��Z4�/Е!���v��У&���k+q��$8��7���v�}�S�؟�VRH� .��j�@����կxW�!��y:Z����Dk���<ǍaO����ܧ�0h�Q�E80���h`�[�����>�Gr7q��$Հ6ӏGw��骮X)I�(�B�s�%9-��q�����kd�T�_�S2 .2p�x+>�Hc����d�u:!�6�f��'	6t9���,<�=&r��L2�;���mH��$I�@B��׃"k��$%�"���s��c���	dUN���S�?W����=�^�5�քy��X5�����M��Du���m�H[iŔ�k| \'��VGL/����`�"ﳠ�|�FY
L@{)�>ׅU��=*����2
t\��K�T�`a�vN�;����
y�*ow�f��J�O�C�j\n�(׆q}��ŗ����E�ė.}=[������>D͏]f�Z��X��x�~�����>�k�����bv^�}�<5�,_���"�TZ\�P����TL�w�5��)�9�R���=jz��77<�Zk�d|�#E]�x+΅n�<��E K��0�'k�紳���>�{�OJnEg%f�u���u��	]%��M�8r�����>�a����F��1�E[�L��ا�O�6�?�� �T�) �(��d��]����V���~({��V������@!,,�6��y�GI�J�E	��=�X�Q�=��\UY�s-�����g��so�
�@8Rx�1�
�N�=9E�A�:���LT�0�0��U^$8I�ꅩ{�L��@�s��tʪ��*����7��|t��p�L�M���4S��)�e�X~��(q&)͊Cc�
j�c�HI�v����'@-ۘ(ʑ��ٚ6���HOnP�=�
�z�*�m�ɶ�&yn���b[?����!�n�,1�Lșa�Lf-n�����߮�+^HnWNu{j�6��v�h�e$վ�h��=̤���K#�b�"O�Ѻ��}3㞄䮭�a}�O���基�NK�z.N�n�ߥ0���Rp��{4By1�D;:����)#���կML���;3g@�\�M��!C���U�̠yE��x���5��VdQ]�|���b���j@����yK_���i(¶k�=%�m�
��+c��=-���l�$�4E[���K�{J��}ld�\���� A}�᭙s������>B��Q�7�$�_&KB�?��;aY�����O����v�c�_�Y�m���U�3y^�@hu� �|5�J�!��� ��D��d����U��Z�G�V�e�L���p�(% _Vޓ?�*U��rV�(��\�Y�6����'X���$�ECg������)��_��{�"�k�rQ~6��tKuJ�	�y��[
4�lXTl��E%M4pGˊ�J�"���c�䔥���;
�l�J"!,�l@d�a'�ԃZÕM��<C���Q�b���hr�-P��'�����a���W��F�D\t*
c��>�����+�/���j���N?�fo2�W@�D�ɭ6H S��u��]U�\4�ľ�$�;����a}T�$]M�A��;;1m���0�&�>#w'�E�3z>^�^�ۼ�1n���6MCͮ�2b'���j(mA^Xv�u(ԉ?C/q���v�-�������Ή�EE�k^&q�좳���Ɵ��Z�3��iW��ʜ��y%�.�o�L����5��sK;e-��SI��r���t�����v<���� �dr�XOu��5H��UF�3L�����H��,�du�78T�@'ţt�Y��f��S���O<�0�6���/�V�.C��5fn�F��]�z�o=N3��Z?�3~�	�R�N��^<ۧ�"L���xLmpX��0^�Mz��!b��K����~m'ۖ�{� �{Vi�ŕCOƒjɼմ6=-s<��rF�!�����^���y#�$�Wʶu_H!oʊJC��ˮ�A�L�5��S0�
�l����g�r4�(�}�ja04e~��ֺ��B��E��.��_�Q�܆�FoE+�XG1��93G�z�M���dB�ۊ��}�d�䨑B����ч�f�ka}ʯ�b�	�Z��O�*���S�+^d]J�ZauN�~���G��g��^���s3��3�e����B;�����tF��8J�h����-�� ���8�?{K8��T�vYdJ�����3��7�h�[	�D���s
��VĮȤ�H(��X4�vJ7�ү�g�4c~���zGL��@�v�����D,�s����j-�6e����(�Pw}0�?�c�LV_3����ݫ�ꝲ?���<9�:Y�.�$�w�^/eq�2�!�N��j�$�B��ݥT�ƪ^8�?@\�E�D�?�ǝ+.��&����
7ط
�aW�6�P!N��#�K�����
WmyX��KHD����,m;�DK���V�=5?����l��P�'�osAt ���+˼G}��!��� 34<�_��Ht�)|���O��':&=A���U�4�1=Y'���,sXZM��|���u�J�-�aS$��c7���7���%vx��f�[������:{JːZ�&*%,̻�́�&>�p�#¹2��MVG(��Dp�v䲰�=���i�̝Q�E�*�R	��;��|��c+_N�W׹��-�*����l�6<���"5Cz��@Ke��j	#�B��'E�(M�+��C#�����/�`�c�$�ٲӪE��<�B��x�_iI,ڀ`�u�
#����/(vē���S1�b�����W~ANUc�����O�VB�In�Z��^�{rOꈒI�����p���
c&=��+Gg&�^��t�n��6�s��S�4g!}�T��)�p.��aK�3Ѵ ��snB�ʛ��)).�F�w.��$=Nއ{�&E!�M�B@���ʸ9j���ĵ�
v�o-�;���U� �I�CF�}�Ш��gq��ڃ�Sy�!GVC�3�|�)[��W��}Z�r�w�������������}d$tM�_��t&JU-�G`*�<�u�SJJe�0��gu"��op!:e����Ϣ��l}k�g�}���e��u�d���)��@�}*�c�����;+\bzz��Y��'��P%�ϱe��~�j/�)��s�ەX�6"����Rq��V��49��K��8P����v��ǟi���ޱl>�JvP���ɧ��j尨-N��Ua��h!�ӝ�n��)���6��!�Mut���U��5�{���_gE��$�����E6�h�N[��D������p%Y�n2�Ѳ��7�'��ѯLַ��	-�i���P�-2E,^�<z�
�F��	a��C�����?=8��A:�d&���k��{��P��]���ē��ko���џ��`�w�͢�����Xshcr��n i[�>\���ҟG�Ia�X�������;����^�l>dc�x^��N��S]���,0���=a'Gͣ�[<������P��[ *t��L83_�@�-FU�Kli����qK�o���t�u��Cm`d���?�eCc-Ttxm]ʚ�g��Xp���������^�����6���y�ml=qk�Z�Y�2�S���ń+6uϊ�#a�͈���~��u��VpK�|�Ώfk<)pk>��gMݟ䤉I���G+�ÞU��q�BQն{2������eI�C��O�@�KK��ey
Gr���\�r�mS2~�Z���~����߯:�H跀f< l�/�{�[�>�:���~qu�W�CY�{��D-G�:��f�Y��-��A}�Q&4��ƀ�,'�]f���J���T�D�&R��;Pha�t�]���ђ�	ΖX0�Jt�!Fa j�fM��>�ɞ�����Nΰ��ѥ����8�I�w�WG$V,��sv�#=�F&m�����$��m/Dݱ��k�x�up���-U�P�l	��BGPt�bd3{�ܱړ��%>QMu&=6�U�e��K���7�DN�;hH���F��Wvt6R�	Q����p>[(h����w���}=2�C����6�T:�� �s�V�'s�4.�n2�M5�832�Y"��29�(wu�a�����p)/���3�Hh�8jCN��dθX*������%�����<����y��!��
(>�M���
�j���~����U��j���ER<(�]���4�X�l���� ���nM�ܱz�����[֠�;U��,��3k�� ?ïR�me��\,D����.���ԉ�}["=�{�@#梹*�E=_ս~�j�\p_;-�H�a�I��I��q�)N�i�<y͍��Y��l�8�?��+�]��5qQ��y��\�r57��*l �x������B��)T4�Y+B�i��21Һ ��O.�Ԟ���V���ߡ�I80�l`���.�]sb!�JN�שB���r!xr��6�J�Z�1|�d����{|�$
nv�!�"{/�8O�rn�bP�M�>>�ჳ_�6��Ş`J�J�s�m���=5-�	����-�?2$�)��(��1[|��/�ke���M�/ޚE�����i��o��j���c���i���ޒh �o���C�ea��y{#��q�nR������z�v��e�e���d6jQ�4q�+����y�Zb^�!��̌�����(��ۺB���)�����}�A��XzK���k`�?9n�˰*��g Dykt�ӟ���ov��ov�5X(c������=b�-K 7-�DM�&���	�{f�8�1��k(	�1I>IŊ!H��sl|�x�6�h7`�p�P'��b��٬򠦇�k�	۟��ݳ�� b6�#;|��HɁ��1��6���^Ĩ���:�wM���٨�G~��|-�����'Ѡ9񭿬�a:�Z����hU�N0��"��	�(U���G�(�o��y��۶�c�f}� #������Y�@���zc����s~��-���;�����$79�d8L�J6�d�)Ƶ��d^���/T�CT�{U�'ԥYgN!4��3���U�59�X�P�7AM'��3)�D]<)5N�FJ�U�wG��5�y�u.���cH�DF�b�_��ү!;�嬌m�,s��9�:Bݾௌt"(%���j�p��M:QK��KXT��@�l��,.�q#�5Wܲ$��G���	a�`j(s�	Z-��D�g�.���碎-��o��.�y:"}]p�a��4T�L�GK�W��cX'pM9���2�S�MWs9r�[��$H�^H8�d��O�]�))h+vsz�᎛�|��F�ڦ�yjJ^�>�B��.^�?�@f�*�
�~��\s;��XʟΏ�/���S(آ�8@��1�!w^�¬��$���C�d`�G9�j�Q�I͕��ъ/����x��+�� MZ�g�9�$*�.��E�	&�27�
�o��d��;�K�
KOU*��$^���k��R�y�~o��^���������T^��0%(�GT`Yu��l~k�u�^���k��g��ly5��9�3�?ld`�r|C��3�E����C??��
9}`ƫ��	������U"��8�1����g�l��й��l(B��^�����4���{r/�oo���%X�Y���W4!$��Wz2-������V�K�V+��o�h�h��)i������$��� X^����<�3L7HFd ���ٲ�R��!0L��h��8=K������v�o9c��S�D����,�W	޻y�bcx�klh�$[Q��_�.v�J�hC<��;���"�S4��#�j���l�Wr��¶݈�C*���fN�]^��w�'�-1
�]��&�ܪJ�߲���y��!T��ƈ���<;�)�i��*C��H��ψR�҉M�]Q�R���[8�oSVR�ŸR��ؓj��~�$P���w�S�� ��Ya)ۤ|?�g��9A��;L���鬊�
2��LN?�r�8T��^�n5>�Wf��x���Y��JP��ٸ�k�roɂ���c�7?dD��k+-n�xw rJ�)?I<Y�Iv3u��q�|I��*�-l"���ڛ4��yakn��+&�}��AC�2�� :�����1M�2��jR�: ]S���VD�3X񚩥�`e�/]K���g��oex�Si����m�^u�hU�
��^��e��)s�-�pw�!.
8�z��I,7���1��>�m���x׃�b���a5�?(���C�=X���S1��Q��h�SH%��w��r'nR.��1-\�oz�0whG��ã6�Ob��qA���=����.�j0Ć��
a�#cf)5����M1v�;���hp]���wu�x�l�A�c��K��N�pD���;���}�d�Cp�xޓ�p�n�r+��`�:�Y�H�����;��73�V��vM�\��H�b����������>g߈�AϫZ�����jۤ��ہ�!m�m��V�Gܾ��i���b�/��6��,��A*_����P��`���ؤ拍a�>$^��/���x���y��n�l��H�c�o3���W�o(IÚX���b�c˰=�TNx]��<5��^����X��;�(+��4 ��Z���N��ۧ���_��O��܈�NL�L��c����EC�D4��,������i[3���D�C���m��ܡ�p'�]49��	���׭MP]�0���um~ͬ!���±&}?���u,p���f�q����r�~�t�D[�[F�W�jw�Gt7�)��_��ٮ\Y����ɬeQ���"<�u��J݆%E�^@����=6�yS�Ԑ���t ��ڜ���6O��<�vF�lv�����ag΢��߈f���p3{Q,x� ��s��7K�ʘqA�:��Mt�
�y�R�p�� D��&�X�(X�Xx���8�����wd�H�ϧ#w�:E�EB��w�9�xo���`�i�B�X�+���q�����-��DVt���y�`Z�%�	���"�!��Bn�'u:��H)���S�PI���;(Ьnj$1!0~���DG��z�q��	��c���Mw�="�2 �U�U	�k��we<��ʗB�7�G��(t���R���x��ħ�S�K�3 ����UW���SC���eۀn�ҧ<���v�⁮�11s�}t���~�o+6�TE[���б�q혨"��#�Q5~�:�7��KN�G�gן��C2R�_����T�IU�\C�R�c��"�؊Y�ļ�.�w��h���@����C��%�����=����#���n &L�5��Z;\E�����Ƒ�4�����l�ѷ?��y��&3��Lݶ�*���G��صk��o�Ҵ�%ǭ�M�U�za ��fA��̕�J��8�}l`�0�1�	�۬,���}�;�b��#؃��L�æ�L�S��f�=$;n���!�k�����O��Ȩ����6���aDƾ��L�oQL���W��ޜ��c<�_\!#��S��1��(��o���n���-B2�d~T|[��R�:� �����M��F��=]Q�i��[�z:f�6)0Rp� EWu�԰����+,��Q��f�_Մ��:)�����˷Ub�Z�$�W`����R��� ���ʙ�����qV	lS�jR��(UT�w��t,��NR�zP��%�i��i������ՄN�ϱ�����i��,,'ʙ���L��g��g��v�T��v���8�� S��>#n㕺la�k���\�XȌ���vֱ��i��盻"��E�1�}����ΰ�����@�7*�M_�CG�|jڗ`Qa^�y��N�OM7�ۓ/��@��8����dM�[g"v�بg��\���-�{Nj�,��N���Tp�/o%�v�e���\�4�a���',�k�ƪ:��k)]:`|��=9��+4O�m��9^�W�h��v�8 �z�>��H4U�����xxX]*'A�?>I2�����cG&1��Yd�)Ϝ��� /	����mn�v�2.E���ykҼ�|���Cob2��	���z{j%��Gqd�ׁ?;(��o�f��G���-\�uA��h�˽ �X��
���}���|$�SW��?P�L�����1˸%��~�FF��[�5Lh�|�V��P�Xo`�[�' }�p��X�TfM[�R���֝S��l�s	�t���`�0i�ɱ�㏑�e�Ⅱz	�Tم�Wy�c�g��`Ҋ��z&�n�T\��z���R�,E���F\=���M5�U�[�����2�U�z��їǼ4�؁K��p�gD�u�5����U�0���R����2P��=��V1��E/�R��mg����v��<�/�s;��]�،6h��K3�+��kE���[:�Z�x�M���ٲ#�x.��BX�dI��[�nq^��r����q��$s~}Ȩ��&/�����}�R��{�.\�铢l��OU��-�E�Y�'`I,�HG��_��d����{/�A�3��Ҳ�6����qDG�J�6��Y@��h��%�����4����l·���b�H�U���Q!	�^�O�c�4������p��/��M��a���5���~��U����|�ə<�����°&�b<�D0	M�SL��U�B�}����r�y�ʯ����]m�ÕUr�m�$��4M�>ä�!���?��2�p����^>��Xuu�*3�@"����e�є8)n=^Gc�/�u�M��u�c��UF)l�57��e=S��:��T bm���l��{0���[V�(�z_��1l����6VV&�_�x�U���(�S��8�k-��A9Ơ�{p5�J�i����饗���氚���!����dV>��u��q��zR�F�JU�0J�D1
���
�xf��6O�pasg��V�?��R�\�;^Xξ��8��u.΃��fi�9��a��&���Ėf�J�\1)���@K�AόJ�W�i05�_@���p������D��� �ު`�Uq���w���E,������>���������	� �)M���[�������	����o�;D[.�%F�Xg���yAl��7Yd�>O�,�D�*�X#Fi��b����#!ϱ�/2L��ޏ��$���`j�ߠ�<��}g�e��A�hay4bgS�;�g�|E�&�v�^a�R5����r3C�hw3��T��5IW�\U�Z)I+�#5�o�D�jq�Mt{m:#}g��o*<������Q\� ����..�d����K裂nQ��Y{M86mQD2�]Џ����w�.�I��������x�[HH�P{4����{o�nZ��w%�WhpŹ��v]O{�Q �b$��Rl�)}A�$���	=�`�c����t� �]�%�.�RȘ�ƫS���Q�	u���x�C���劄�dT��J5�0Ҟ7����u�1�����5�;)�=G����&s��?�.g#�����H�.HS���k���oJkg�ra`N���Y�;�N���7��P�g>士�LP�3@G9[>g�7n��V&/�ۮ��&[OwA��S�wʱ���O���a�\5�3��Q.M�_A������f;�av�w��
8�t�;3Q��OJ�:�A�P��6ڼ�&�h��iW!©�Ζ�3�������R@+Y=�'Ñ�刹9�m`��X��d���0(p���\|t5����S��u@�K"��#�3m��3^L�ƛD6TaK���9��H�N���,���W`������	�7^�ѱ�!��]L�?+7��&�ltq :ˈ%_�	7���Gđ��"_؟�"�G�<!�/����#~p�B�����aWϕ��t{4#^PnYA+Kw����O��VY-�a�;We{:r��0��3�%C�����{a�*r��x�CZ����mOz���4}JN��-D�CM̤y�n�g���r�Zg-lu|��O�/��g�K/��Kbل�vv?�������̹y%a����)*��6]Ct*w� L�����{x��/�abGzb�E���p�չ�B36�p�sxRޫs�<#�l�=����s~]C�q>U�!���yLu9)����� ˫��9�~����g Ե��SHaZ�ǭ�HQ9�4;�ջ�+���6����{W�C&�}�YΦ�i[���0��E[O���?�Tld�gE�1�;+5LW���
����m��J��&�P�1�Y��~���!�����݀^ �T[�-�>z���D����1����TL<ګas� 	�ܫ����%����x5(җ��*��@�%B��&����f b���BH�� ��;KH��"Ǯ�F:�Eq��^w������NzoV�>	�A	�f1r�参���8n �� �W_/0
���w[Qs��q��{��O1|�{�٪$��3J<`���������6�{;[$~k��L�y4����fH��*f���V /E;h��*��~��]��PW\�#}SDf���Q�#=�}E9�������$�֌ /�ڙ�a��z�.y����d�2A���~c�G6C�ƫ�E:NI(�ź�-���8�%Ғ/�r3���R�R��32GC�����aZ��}�꧅ʘ's7讀�V�s�J� &a���#�o���.l`�D�����uӹ�?
di�E��ɲ%����$��m���q~��ol"o� Y�WUn����h��P��9O���\�����/�8�߽�yOn���;�#E����Tއ��Y�$r	>W���r�(�״��vU'����>�#a�f�l�4�1��y��Uct$~|蘴4?��r�]0yZ���v��P��0h��^=�2���98#1 R���?v�9/��p:�r���4����L���h�IrU���{_j�a�
��0~D���[fR
������l�r����֦�e��C��{��Y".�iO�����2��k�Kr�Ӟ��_H،���x]���8�M�`4�%;3.Z��g��~X4m��2_Um߄�2�
�&��O� D�X6��Ǭ,�����8
�M ��N���+���B*�\��R��;vWR�L�u�g�$	���{W�6�p{����Vu�䴣�bA�j6tm�!����S5O�W�iD�Ae�B�U�酞C?7*�f�O�|3��K�>'���B4��q;-�\nx�WM{ ���Z��tT�V��$�UI��<R@����o���.�G�E��>�h����a�(��|�ZZs؁�),G2�,c���LC)�n��	�92���6Z��ǳW�|�=��	���b��%��Ԋ�m��tGB���i�y���������6�P��[F���{c�dYhrt�k+���,�8�ľdzȶ�h��0�� ����\~��1L?�0��Ym`	T�y.���n�D�Ǖ�R,�}��jN�)���t�͂>E�0�Zr���M����za��-+NTs���0�K��"]����;��|��G���^���具�ID�v�m�2ְ@�@۰9������>a�'�\�0%��_��,�s(�zu0	��)�	�"���-���.����S��|;���6���1i[t�<o|h]6�ѵ\`&Y� lXN휼�.%� ��5df����-�<̉���ޣ�)��踩��/E_ ���d�������^��nz�F�z��.,�U�	WHT��!.��2��*��
~����l���'�GE�
���װ�f��Dj�s����S��Dg$�m^�҅Z�(��f�����z��x�	��k]���J�*6F��}"��
���Q3*Q���"�=�O$�C�a^Ή�����7EQކǐ����8�����E�	�o ���S��3ec23vP� g�Q���H\U�+���u@�>ی��:�V��ʉCl��Sr�AE6��Zg`;e��Zt�<�|ɰ�;o�[hT�.�*N�I����ޙd=#ڻ���)|*
�_{&�T�߳�S��vj{�|��f0�
1�o-7�c0fp��)��1\Sv7�M����W�)��*2}�l<u���a ���SO�~�_gi�I0ҙk,3V�҃]��d�C.Qz�rW��楒O����#�u@�'�w������=��`��9d��j���y����vBIh�`LG�J�{��e��< Ŧ>24�/}2�����/��t�r�����"��g�Pcb�8%�i�l��)mN�>a�������h���?�6�S�s9/1����v�|x����ߏ'n��`U�d�Cb���<#Lv���%d���f�㥄���N�����n��,�Eg�Ȋ ���:5bd�غV:�'�������*bh�d��R�T�'��GV;�F�!�?���c�	y�,@�-:*�s�E��&=����9�n5':	���l��6f�-\��������oډ{������?N((b"�,���'��X�d�tm�D�MT-,0�X&;y�G�BKs��'��h��]��T8�Z�I�x��r�O͘�t��&ʘ�h��w�hF�����u�Ow�V]�mԘo�Q�+�PHTC��϶��B�Tg>P�p��ߧ�h�ϴ�rW������tU�{`>'�ҧ�CA�v�9[��u�<��[��OQ���#��;)�j�hi�b$�ѐ����Y����`B�Dw�A�-颔N�����š��gO���y�5�Ę�`6��D3�F8+�ťqSi ���.{�u����_gF۔�-���Hc@:i\3]�Q��}S�\��l������<���1[�E�{�|ʵ�-�8����,vz�wٴ�`nj������gЃ���=,JkWC�����?�4�v��e�`�ɴ��:��$#��i�8�z�'�ʫ{�;{�*���r���@E��=5\#�AL�,-j^3�S��T�	E]��EL�6�׀)��_�\���!`�J�0�d���#AP�K��A���ǩaC��?��Ҡl
���%
3�%Q��[k�s�a��ª��k�	h7������>'��wE�=(�
��"K��_�N�d<J������*
� Q�|�$^���ky������ݤ8�c" 1I"I���_��q���e5oE(�<n�=�ڔ�]B����F�q;�&��Z���}F�2$�2]�9Y�E�Z�4���Q:�6��*:ک-e�p)("� �l�s[)񲩳�\�]Ǣ�X��ߨT�me�M/�*���*��y�T"�h�����r<�٨�~��T��r�&̽qIY���0R����� �/F	טq�J�
�4����Y�X��	������29x�6xgk	q5�n ��R� R�!�
]�_�G��5�pFn��\ש����4 /�-DM��楗�RDl�U��{{g7�V"r�k.�c�����kƁ��.�w�u'Ȋ�oo'��C�s��H,�-�0� RAn�r��je9���H���]6sY�xz����W��(W V�4��4[j彵@�pLU5�r�DOZ�GB|�Gp��xD����y;���9.��U�u�X(�mr�����X})��'͐ڈ*�ǽ()�?� V%�0�"vf��lL�`�zK�<���O�~I�>������(��p��Uv'ZW�$���Q���{"����i�,���\������j
�2A ���4ا����JHB1��*"\����h%�-��{{Z�D�6�#ZÑzA݂�nV�T%���x�Wq����tZ9k�{��[�����	"�0��.<U �	wgC�Fu�a��"�D�B�7�-�؇1��~�w>���xV����C��T-sȏ8��<(Ʈ y����w�$�~��xñ�2�ńx��[)��i��H�x�<�;1�y�{!�YL�*�,4�cZ;�3mkޭ���~��G7P�XJ�QQ d!o~-���P�Yg��F[��<?w0	y��%�I�ZZ��% �~�����%1�hO�a���S
�"<ܢdG<���X�1ݿ�ډU�6�>�Sk{�o������ux�����Z#�t\�{0�G(�%�~%'xi\�x�f�`]k�a��� ¥��S}<֦�o��\^p�`��f%\���|M�a����R�Aq	O6X\�FZ�=��mƯ,��މs��]"�D�B@h�!3_NB��`�l���h'`�MgC:!�)��?�u`S�5[�uF�p��!e$�?N��\D�y�2gp�o��=O��QF@�b���Xܓ�_���c�6�ފ���e%�(�B�I�ܝ��f1QC�%NV�P���(�G���~M��OO|�������_/�F�ǫ��@��#����H��v�@�I�v#Z�.?V^	x5w�H,SE�M�O�R�wbh��8&�?"`�\��6�H���cq��kZ/I�U-����
~?4��V����Ri�� �Z�����#8�$�݊22̶�jK���һ`����lbM
T4WR����ւ�aGBKy4A�|�k]*�r���Qr��	6S@��(�gс#c�oc��o��]��uK���8�t�1�<lc��H�i�dW`��Go<�1q%�\J/E�Mi�v��Y��\ʿc-����"noP�8�o&i�	%��-;��.���b�'���ݹ�/��N:��@T&[+�������t�3�n��xM����ҽ�v%`�gƈ��I������)��ŏ>Z	{�8��n�R�tZk�����O`�Qh���)F2Z�=Ϳ���i9���4w��9z���p��R��?��z��a�.�일��紤�������u{�C�sB>��4���*�z��2�)y�~�ў*Mm�0��������r��bv����WwQ�S��N}톙��:nl܉�Brˆ5 Q���(l���/P�ޭ��9w�c;���y�$�)��쪎�H�vP��F�R��e��O�����G¯��S��Ƃ� ��h��Y���U+��Ycn�(L����@�}�A*G�vJ�z��˶5M�,5��h�W�Hā�����G�Y*�)x��P�Y�l;#mN�IO���+k]=y�W�R�b�h���c
�eW�'?��5𴧗M��������f��!��i\8ʦ��7�eD��26�A��ً�\3!"�T��M���+O�c'15�������2��n��^����/4FL'?YSL��jb�w?�X��(��6��Ģ��M	2RV���G��0sÝ�|���&��9ZP��%r�a��G*(j�i���a���Cd�֭K>�ypq_��u���G��]f�R�۬���I���D��u��Ţ��D�5X����x�Ɍ1J��ƻ:�+�4���"sXgfH~�����!���W(L��aL�.��ѧ�|^�U=�s��������8������Q�u����w6�!"FjpԲ��l�l�a�s�U��g�H�H�lw,�G�p���d8��l~�_c9�M�4�dV
�z%���1��L�u�R�
|�G97/�sЖ�_��OTk�� ����S�rAOO�B�r���e��Ƌmx���Sٵ�D[�a�}�0vm��ؿ1U�5�b�㩫�4%
U�Cګ��L��K�(����V]�5�Ґ�I��{[�v3*S��Jyku	+Sȿ����Ծ�%v�p7����)&e�b����(�-�<�R�c����,�{��UNQB];�,1�ϴ'�m+�896"_R>��#=�[rd3A'>�����X����'�޸���Y`e O�yh���?~�O�+���ą��u}� �l��@x�ae�'��8�7ڣU�N_�&J.�=�s�bl�=�����!��Z��@R:�j1"�YU�k/��c�E:�7�g/�K�8�#:l�KH��Ϋ~(6˘;ɝ�D59�b�o�nP���/��qR�qS�37� �N*�"naQ�s��6I��ݧx�K�?��BЀ�2��5<���-�(�3ߖ4F̶�ȹT��֩k��t����J��b�G���� �v�;:c�HI:n�\b(1���è!��۫zP���K�X;�Ѱ�7x�\ܾԫ�j��=/$��e�)z�����d�]�)����HV��<b�7'���ܢ��*��}|Gb���D����ky��'y�
������{�Oetj(�	\j�o������b�Q���\�N�yD��uu�}�~kx�bh���a�1$
�c:�9�vZ�V����C��?�Np;x��ˇ����[�X�����~�f�c�~&��2����r WQ�('�U���ωmX}ke5�|>�5���+pF���%��O�"���#����?4�Ҙ�������B��!,��������!Q�@�v�̰��]E������gc���;֏|N<���w���^�J���D���l���pfK��M0ؐ~�Շ�{843�w�_�����jB��P�*裌�G��|WP�����?�eK�)6Ek�L�J,�Ο"O��%G?�m��kX����������D����������]qM�F��ۨF�yN\�7��rH��e~"RXh�~3���I�[�"rL�Cd�l�.�F�5)�G��1v�"�9�sbKQ'���KDM*�
�U�+%,u+C�f�Qs��@H���/9��}�*yc)�:7ؚ���b,�ӓ�L���՛�V�y\��7�ry�Ү��Jq���맘�E�t�����h�Hho�%�b��n���+��H*��5����B���lWy?�@��D������ȽQI$gĳd7��_Z;UU�m���k�W�d���uǋ�|��
_[צ�%�.��cv�d�l�� �F�[{��� ��n?2j�����)y��>qgVo|�;� ���8eI��.uhKz���,�'}Q̳t�"	�=�;FcA�h�*��s���b��~�%�LӏgS� ~K��O3s�< ��jd�����
7	)�V��s�v�����Sh�.r���N�d~�r4���́O��dr�_�9U3BB�x� Rn��O�1��1�<L����h
�J뱲Ct+��~+!�%�K�ּ6�&ə/��7q�U)�ҿh��N8�3�촴��YNԢ��E	X!]~�z_��^8������`��o��e~���f�������M�m}NR������V@��{���e��TN��������a^�y�����N��L6���w[��ޠG�����9�9e�����#�K�!�\�[�V�P'��z5�h
�ˍ4��ĳ�!Kl�>8/��G Z���5��D���������;��ɔ`���U��bf�aV���P��.�/yv킥kߝ���q��@�70��,H(-D����
�/o���MӬ�b��zk���6�>9z��	����֏��t8O��Σ�g��?�H���u�罯��"�fT.���X�R$� �W��"�g�|h��(P������+I�(6�����<1-��Gm�J���4Z[��]x��U��(:���H�e±�^��wq�hN�;\�p�׿ugM�}��Q�o�+����C\n9����&�[��}`�xfa	a�����G��Kz��:����ӥ0�,2��L��k�&�Z>L��� &��[�܏ {��r4��Z3��g�*�K���T�82v��KPc�
�̈́7<]��6,��ɈgR�22�w��~�_�PxG�߂J�6q�J�!|���l�=z���ڞ�ˁ=�ĐϢ�0k0�n\�Cj�,?��!�jT��(���'O� �R�� фġ�T�T����ʳ�[ �̩{��K��ڶD�Y8�l�r˒�"��o�(����*9���2U׆� ���#ψ�9�2�*�`H�s�$c�,���VRI�+��Ϫު��>:���=�O�%�lΠY�2�ș���sO���2���Eֿ��k���Gm�� �y�ʹ��j]f	y��<�g��z��j�T��ԙ�ǃN� ,�TdB��,���UDi�I��V���o�6P�@P�٧~���	Yn�D����XV�ln$:�qٿ8U'Ӽ�XUD�Je��Hi�>�fa�G)�Z����f�ۑ�,;���u��^S��U谘V�'�|I�t8`�p��t	
F����D��4`,'�T��C��Õ�����9�|��h�+������:��l�I�tN�a'{zj'��±0�> ��O7~�U��{Z8���n�|ԫ7�0T��˓mè�����H(Ln#��S7�%�&�� j�w�.T�PXA�~�C�_�c���f���.%�9u�e�c�����Z�ʑ�_6��q
Xr7��p�m��C���Qs|���X�@�eჁ����Q#"]c8g_<L��2���N_!*[U��m�u��2w�*u�����m�E,�
��|�qZ'��+8��KT㢄6�\���cR_L�G��j]��+0��(Q	ڨ����X���y�D�!fQe�k�P$y�7#�LoI��a��Knj�u*b�~{���L�l�=;esI8��e6�i3;cᖖZӊC,1�'�n�Y����B'�7c�ѫ*.S>L-gt�y� ={���=�@#d
]��&l����57�O\�m��3��w��-F�1l��c6�Ө�o���e��&�C9�r�U�	�N6�2���ɦ���dȀ�E�u}�?BB��w��H��NM�n�֖.ؚ�3�O�"ьB��A&���첒��N�Թ����_Q�Ovw\82ޡa�y#h<�9b����O�g��^i{rE�8���>�b�\�1�5:��:���F}�G6��\[��f{�anko�8B�3�bO��B*Zu�e�R]o{ҁl�D�6,s�P�	�A�G�G��
.^�3��(2I?���椞N���b�ĥ��!��~�	�����f)u�2���	�F����C:�8E��}�Yg��[u-�2(�]�M�\/�w�X��+x�4�K��
�阎~d� ��'��Eo�L��j/+�r@��^,oަ��~����UEmI!Od:��sV�������-5�k�����L���� ��aK����%t�i]���=Q����-�8�wu �Y�S&@�9�,��u��f����;�d���ʼ*@�l�j�U���3ED��j����]v�;���Z�=�DQU֗�#�¶j\Ι�,(��G�Jy�dD�.�ҋ�-5�S�}�r,�Č1ɭ#���l��wh5�Aä�E����.��hlYW S����sGc���`�뀄�W��t�5]�%���	��.��0v%�?�?l���=>̙�0G��v��E�4�0��fV��M`&��xQ�����/����0�)��:�ԑK�q�1��1[��"��b�L�D�D*�AӜX�yDx��i�
w�>�&�z
���S�M��ÒQ\˳n2i��������X�z��7������c�������� ��P��6�H��X�pT2�����s�u�f�x�)�͋/(
7-�L^�t����ݼPMz�jcDt�� CLA[;\욐.��3&"R\=\���0 8���<��X2���_��J6��©��ҵ=-1k'IZs籤�\���n�s�|�g�c�}�c�#�CH�u��Բ�}�y�^�P���fN��&L��O��`(	���h�[����3�`��{��7t���'�r(��ײ�첈�{618���>g?��`�XDWe/4���JgX�aECX �_�+I8'	vi���� Z(I ��;��Ռ"9�I��P^� f0
e@ pU�����N�]��D��Մ������j�� �z��(�J�u��ﳠ�����A��SX7+6����,f�5��{���00Q�]���y��>�r�V�#� �ҌJ5�p�g��s�X��4�&��Fw���C���|�ـE�!�y��`��L�8Qߊ5��z��W!��e�W"��6���U�<7���� js.�{=���_�>/������!'"�4�Q�̩����#�s��Mo�}苁�Z4�f�q�Ƨ�P�i/�����<�1$U#z�sGh�S�:��cl�.��CXl��F�����>��C;�ҙ�~!xzSO�h�u,EV.^ź��B�I^;��3x���l�
" �ΐ;��8Oxm�`�b<�X8K
�:�Z�&ń���66���?�:�H+�5�n1<���4�2�4Ƈ[�͉-[e��n��h݂ä�r%:��e������b��J���o��3^V�w���(bI�&�Z�s�17��v�;����}��/��|֨����j��h_ք�Pf��R�y�mb6 �lr�ۏ�r��ōĞ�"��ؼ_,��DN-U����.v��B4UN������/k�@��`Y2*��¯�̬Е���߬P#е����'� �Mt��?�7��Yl
Bw��Mr�6��6�-��<=���O�U��k����w�a���N%� Ly�~�ر��Em
�,E�Ű�[k�\:�0��}�e��)i��s�Z��)�޳Xͣ�HQ��њBL�eh��	I��� raoH�:���g��Zc��U�I�+�E���Y%n�zM��@Y{�CO�G�d�&id������R�c��J��m�蔊Pg+Zm�~U�"y��d+g��:�5�~YM�y��f)K��;r�]��B%��?�4����x��YF� 7��kP>&�e=��ՠ�?"��z��q�３�hB;}����#�.`�C��(�}�T`����Y�CQm[U-��o�|��ev��vU�S����,�)�%��2Z=���6�O�o@;t-b��m<j�II�~���ˈ[Ggn�����t��O�J`^w9����q�ԃ���7y��e����e_f2c�F^7�c$�&��Yk�w2`N��n�E�$�Kr��/w\?3�
��ݙ��Du��ߏ�v����\߉5&����p�������<L
f �0��6_I��]~l2W�Ќ���>,BF�5�b�5�%,����bU�ҋ��
��[z�k�$��qV6X�b�3Yz,�Qm;�}Y
�{5������ad�AHɝ��}��txL�6����|�\����^zm������̒^���:9P�ORՍ$��i'�$��[�����4Z`�6�;���
c��[�Y5��RuJ��q�(7Zm���}���+n|��&_x'"� ���;×)M�P�$� =س�4Մ��O���7i���|��DL��;M�rmg�ul��<	plK�k`�k=�=���C��� ����	&�0R�F�P�Y�<�x�� {4�v�[B�.�����tJ+�t ����
]+�ÏP��5
���J�N��^��&2k���[�Ê}�������˾���sPP�Z&*tH7�e�'�iF44�׫���N�g��9�EL�8��Qw=VClTO�d$�
�Ȍ5��,}���)��5��B}E+N�`6��/�W���UX�j�g�w�U4�5r�btf���~W�s��������Z�xb�L�pB�=� �u=���� ���Wn�f�]�FǛ*������6�@���CV6ޡ#�.o����]d^1��u�
}�����p\i���L�mm�o=�LX�	@Ч%$�m�qqV�_�'���>KX�@H��8�<'F�(��R8"2�E��P�nT׸ 0L�/��Qu����NQg:Up�fT�[��γ4R<L���T�A�:�hK�St�t����,�\2�A��S�h�E��'9�������$$������ Ϩ�r�:��j�6�� y���ޑ����6��jI����G�%��L0�wI�=�1ʁ��Ұ8j���N6]tK�.��i:鴣���鐪�j�XZV2ْ�mMh�4�x�)�rZ;�~`�e8N*���#�4h���k���ѕ-2��%��ӝ[���pn��}�\��Zk$��E�I�Æ�m4�����-Ib�.$�c��9訫�h&	,P�x�U�W��G���kH�lhw����lJ:��V) <�hA�Y�س'>#Nk��N�&S�<<�~�]�eB���Wn��A}�x_6�%V��{��-vJ��M��-�uk��K��ޖ��`A�*ĳ�Z;�Qa3�/�紱?3��#Y:X�?Y��0�k�8�_���4&mj�:@ ��v��\���b��*5�NA#9���ф�V�4$-h}�)�îڽ�O�$5t'@�$�R��Ύ�X�qb�B�>�����%٦f5I�T��
A�1B�MC�;P(h�at
H���O(R�V�"����;�r�k�������Pf>���P�9s���?%q��2m����ZMl�U�{mw������A�7#�M��Ԟ�S\��Ю���F�}�F_���6ӣ�z���f�L=�̃�EB�O�!Bj+qN�yc�M\x�ŀ依-~tM9�6vy{�7�k?v)	���{��6� @}�F�y�p�ދ,��GT��Q����>���8���c$�Z|�O1�R-�м�цl���^����ޮK���k�>��ѯ|�~���^�:�c֓0oȈ'�+2\p��,ʳ<��|��B sA3�g"-M�zy,��:e7/��}ѣ?D-I�KvWɒ����u�
s�(o��U�	��P��]g;� hL%}Z��Y� ��SIC�|�{ezs�m�W}<Gl��ؒe;�o�"#��u����%��ݎq�A�d	�uK��}�������A�H�%��u}��uް�B��T��'o�� Xw���!r[NAAv����xu�-�����c�d�<����[��o߿qra���V�B����Q�U�]h��${���X��+|$�u�@��ܧ�/ӿ�����1/�6b+X����c��i1�Hӟ�9'6?�Ě٠�l��|û"��1���}�-$̹�!�NL椛����"*'��Z֤��_�F(L�%�[��o�V:C��$,ώ3f��}�߬�34�E��B)�V>��:��=��{
 P�v��z�2u7+V�=\𿌜������P���<�	�������V�y��m}G�?q8M����0I�K�Y��@�
��uU^Q�FI��&,�y�뾡鈹��Ɉ�8T-1\9i����2r���*/4�C��p]y?+��R�	4<L��ͧ��^��Pb�^09��X��?��qd��%�����[?��sL�>c=�:Rj;u���&��E,�M�U���n�P��̆y��gp	�h���P��iƙX�W]\�n��QR�j���I ���n��$K��I{���3�\CS A6��ϡ���	�Z�j 4�LZ��ɬa��0D�\+��J��i�"��Ɇ.8-��7�s����e6�,�#��lJ����̀��ij/&K����<�&�N2N=�5�&��{i��q�saEX|`�V��&�n�{�G%��*�?G�T��d�h�[ ׶J�&�Ŭ�$X���2tʧe�z�[o�;T�G�5����̋����ҷ1d�{�7�B��ѳ^O�[�)�A�1��&��rtr��x�U<�����*��W�-�r���6T;����9�ޘ��F�k��k�À�=f1���/�b��x�0�=:U�����[��4�����O/�*�0N���[��� ͥ�mY�ȃb�!�"ȭ���6Ƣ\���ԣ(�8	O�%<y�Bt��z�V�Ur �6?oP����k�NDIQ������a2�i��}� O��aO�����fA���	PF�����Fqz;�`�g��ղ��|b�H��j��#�N@K��L8�~s��e�fv Ȕ�t3�<��䱑BJ�#ˎ"����O������}Н��X�x_V���\l�g�"��ڽf�}���lhIz��Z��%!D7B���x��<x�@���e��y�fR��ٲt2��-��+�%ZW]��[�:��f�+�!\�ek<tF'�1P'�oHg���h�ƌ��8"G��M�]y�Gm�bv2����&9��W�ܵ�cS���������c
�6I2��[������lcED�������&1�����8C�jh�gމ"�$|�e�U��k|��^�Yv?�`�T�OK�_�x�"�$P>�#D��n{���e8_�d�q6PFn�j61�>�sw� ��cZ�M�'h���g� ��_��ZTOK�w_�!?{������F'A�@~aDVĖS0SF����G>�w��6��X�=I�6ecJ9��:�x͎��ڢ4<��W`���7^pC�_�� $����!d�7�*��=YF���m�ی��lkLֈ��Kf��H��iV�畋W��pD�}l&��'���p݆S�&N>�$F�g>��!�˟��S���q��C�P���qp��M�xl@	��=��f�ϙY�(��L�ȫ��Cu[�]����h�	�6��0��+����o�2��[!NH.Y��n�a�8�v�E;�y�t�kS_(ӕ�Ak`�/�'�`m ��}2��N�D�\��fi�)0fP��\:+wkgm����1�G�0;A�,/��\�m>�\<r:c�l�)O�������\`�WTk��Q�&LD0� ������[[9���<��qb1���[��=�{;��B�����T1��	�R��={o�1Z���B"pʤ׫�#Ϲ��
-�z���]f�d��# �y{qv��]����f<ӈ��,l�oA��aj��G�*�1�D��H��^N{ո�R����]T���5�&�0?qg��"�z���KdQŵ��*����N�}d#�2�ɓ�c�s��]Oࣉ(=@-��[��~KP��?0����	��UF�D�hK��W�~_��ܑ��Tͷ��H7��t���ƛs��BEe��^ �F�M ��b_��[�&C:��E&�	{MCv��D.��;
�G{�ů��r���*�a��W���bUa���A����FY���Dы"̢#X����-]�P��^{���Q����}�! ��mx]�*�ҺB�$�YM�E������~h#ڷִ	0E�1���	�۵�A�*+.��q��w��T�dK��q�[�������{���Jaſ@O��ʚ�d�+��W���)��I?��Ư�1�0�ˉ�Q�ё�.k��/���^��0_&]�K���%4��w�.��t`2b2��W �����U>�zVGz���s��\����f]�e� ���ݡg�-�\�NM|��QX&�^S$7C��K<[&؂��;�җih��0 �R�#��d�X�S��8�l�>���^����~۵�������)�a������8�~̌!O/?Ip��!~�:��k먕�¹���b]��v�6�v}�C��:9�m1���9�}��]�t�F�jƴ�y���>�I@��6R�+�U|ǭ�����øxJ�~�NË�`�s37�� Qڒ��ofYQ�q��ݣ�����~�-ro�#�8���gq�j��ìnZ9w�L��X����p�聦.�8�H�F�+�6*!56�A	[���T1�B4�M�4)���g��X�����1 ��M��YbcfbM.q�#���̘�=����A���TjҼ�ec�IJ�;)�F���8�Vke�ޓ��� �	��p��j��Sq����4I�P��
��j�m��L� ��X��A�#���D��웵е#|�
J=
�v1:4]�2l���Q�OB�J�;��pB��"��%8�s��`zE���� ߹����h���+''�ex@t$l/��DV����81�7�5d�����\Ա�q��q�e���ܯ$���d ����{�4��^E)��Ys�*�4���߿�93�۴�(V���k%�D2�$H�̚��?H� n���U�k�<�7w
��Oh�R0F͊�Tb��+��ܻי��.���b@ٙ���+7�jp�?v8M��<v���N��F���!0�$Wp�� x��r�� �M��x+��X<�V32��3�2����t�B���Ҝ�}k[��j뚱=&~�
.**`��7ڏIr��R0HLXl��O��� @݌�l�qK����{��;k}ʥ�wm�8�Y٧�M��Ǣ�Юh/B
�ۯRR�2�+��P>'l�2"��(�-��^�Ap�u��>i<��
+��3O7g��0���h�1V*��
����ߛ�s�g�|�dV����Vwϕ��'��u��8S	��`1��M�o�� �m���g���#D���Om���)��QA�ɖ�䂼qb���i`��_��<)�L�<���H�q�r4U�O�o�����1+�gh���@�w8E��I�Cv��`=saZ������T'�z��'
*{hH� �3B��h��Bg]΁(�L5cǍJ�~�i��H���?��c>Γ�)AgR�|��^��.��C�u�������Ź����s��3u�G&�OL���@��O R���y��E��vRm�ih�]�'�ı���[����X�5k㥅�P��A��@E>�}|0HH���_dl��H���cs��i��zǇ�>i!Fx �CH� ��w�۟`��r���{�|c��Mt�aVM6Fs�QS���C�� �DHhz�Gt��it���hj�nl�dVqT���&t}MtO+�i�5.�Θ�vQ��V:.�j5�
6�\M$,� T}���b�Oc�:R�gL}�:�~��{���ZY��Uθl�}����gC�&�{2��e���mJ'�+O:�i�.�_>D��]-��$|D�8s���)@��([��!�h�d��xjT������wJ���SM�T�&($n�X7������jtD��Ӈ5瑇�ES�^�v`�Q*P�#5�%-W���ۼ��H%^���5
h������clҀL�p'Cǁ?�D�I����s)O#��!��>*#����_�����K�\
̤�Gn����?�c���L��z�W�$睽sb�O��f�^��z���G��,��z��2��3y�lh��^��[���v�#�)�1lI����M�~W^�_1	&p�]�#����Xk���jr��݀�(�d@]r<h�|�R�ĲL�`���#����ǥ��:'�:�k�F�&F���Dn'�j�4V|p����
l��G����e'�t�v�;+3Ϙ{'?P1�1�\��T8�\A�\?^���
�y��}*p��5Ik��]��QJz&�3Ǒ��E����c�5���5���V9��1�y���� b�����弱̬ѩ�����3�)�ӓ�^!�r�&=�t�c'�XCo%���C���;�Ξ�^�ٝѢ�_�]���G+>
��'�+z�
��{>�b����1�.���QZ����NME�7��,9W���p^_�8�]�B&�ַ1.p�����T��D��4^�����Uq�Z�]p�`t)��6i5.��+�V6�H-V�8x���k�2 V���A8�汵�DfBv�]�,�k$��V�#o�{���{�
!���	ֲg!�&���,,������b�/�2�g��<��eFU��=�J~�-��r�BL���$��.o��M5v�6s���NIZ�1a�fiئ2�îm�i���-��{��Y�'�F8i�V��儞3�"���H�<L��j��-d��ڟ�2�������{yhCDhf�*CJ�W�SB������R�}:u6Rp�9eJ�A���TKo��}f6|s����]���0fڧ�n�� E��T��t�Y���#�?c����>>�"�	��9�r�b�7�ğ�ݚ��bzt|�1V�wf��G'��9�Mc�6�`���O�6�݋T���
�BJ�ܒ7�^
�?;%�$����}�*�M3��s[�S��гb��(P�z���a�L�~:���`���&��\�S��\,��L�Y��bb�.�X	���h�7����;&���qĀv�J�����z�����[9L�%��L��k�o[h���8ZԢA�.��8��H�(\dg0���,}�*d~�M[�J�(��.{�kIl�n=}�Л �d�ˢ�1���"ס�Gl�r�w��K��PMZ�8�Y���,���pЖ?�m|�*��L�H�`�Ś�-��@I�y��,��������4���nn-s��L
���������0��ī��%mRdk�ˁ[�©�̀5o��G<m�U�����)Z�D~��j�d1oܗ���<و�`���]�,4��tm�M7r���GAX�6lި�JA��/\�*l2MH�[�nƁnFbt3�i5���Rz>��2����� Ԍ�y�ٲ��������^~7 ·as��u��uƬyi�Ld�����3��9o���������S�.��%�@9�Oq���bU���}��ꑝ��+?��l84�N�N���yj�&��槽|,L���x���֓��ƕ�䥱�S�8�� D�Up .��e�S�S�Hg����~my���P�E�Pz�QU�'igM�F�ۖ�L��B��^��59G8׽%�W��[ 7�k�F��PM���/�朚sz?N��3�5zN��Jn����X\q����K���2u>By�(��!xo��j�#��T|
�=<�r�r	\��o`� ��_����RF�������7R��\/����W��IJV��К���l��K��"��J_]M��M7�)�f;��d?i�%a }���A�W�����{��BKV��m;\�"�;n�ږ���T�=}M�o�u4b�G����RN�����'�����Ϥǉ�}s�@jM�FO�&���������B�)+���8��1����#:���e��xs�1��I����"�驸@ޫ�E1ɢ��`�ꯐ@���6ί[X���Ԑ	 �[�
M�bC�Տ�t�W�c�rEb�� ��O��A�P����s���� ��}�ƥ/���1=�#>�@ӴЕ�����fY/�B=�{�@�g���[(������<�8��$�]1�m�k���63�Y|~��gj�hv�Io�,xk<c
��T�^�]�U �����l����V3��1�Q��AXd@!� S�7��1nQNV����ũ؝��I�p�xW�ٌ	�H�p��y�y���d	����:�������ϹP]��������	f���;��@��3�w�j�W�Q��$G�gxU�m�lx��p�H���j�Ӆ ��a<���&��W����멊=�v��R���+K$�+��淭��˵��u1���{�����q���{e��@�������6�ǥ�(X<`��ޝ�]~az���|&/멬!�06u^�ҵ��m�����gL#�/q1���w��)z�b��ޭ��V{������0ߠM��'"��u!dF��{��%��Jy^�'�A�5���3L��2���ӹ�v=���A���V�����'H8{��N#э|��񸗠K�s���3砩�h�1�o߁���c[;ڈ,*;�OH����U���+�c��0제��7�����4�ٲ��=p8<�<NlWEe�)�Ue�h��f0҈F�����g=��qM�eD�Jc�.\g}��W�����)Pt򮀺��3�}.-�#��j*C�	�����Zײ�&x��$�7ˬQ*LtV B��B�#�5����K��:�@��
�)�[h�k�j�n��J��v�O
�������4���d��$Y��.�3`�f0[�������NgkM��`d� ����v��q��G"ё����	w����f�Q�mp�B�n��� f�px�n��r��))w�J�?���`���h�vXР�@�������m��/7�� ���)J3H���ڠ����/s+S�x6��lܮ��wc3��86��a���'�q)�����j�E"R�tl���?�/}�m�D��3�}|���}�<Di+*�'D�����p�!#U_�9�ޙ��D5=iIJ`w��51�6��3���ٖj��诿:h�vP`�r�����M��_�O�����&G19`ى������]��]s��h�M��<�Պ`\�i�8B�CA��Q���6ǇCG�OL�"���-�d�p��]��-S��.%R*�����_Aw�
}^��Y�lrg�����U(��O� �d�=�m�j,�\cq�<�{8�!L��B��쾟�exM}1T��
�ɺ��9���Fz<O���i�z�袊g���цm�7��FA��Ё��GN�
2����;%v�g	��l���Pv=�5�>
�z�[N(�R,6��4�2���}�\���I���!L����#�v��z�EÖWr��
�Z՛'0�	`	0k�=��#:gt�b��~&BF�Osb9+�!I�������Mq)	����GvQL����<��Y���g�W;���KJ�7v��ߣvj���@��hc��*��ӈL�JW�1�/'�2��'zSF�	 ��O.��qR�,ETQ?�ܽTz�S斜������1/:�"m�gY_�����@�1�/�X�ҹ�4XE�<N���D���̌f�E����i��P�J������Br�:�s8�Ҿ�hj
Pp�y$���^^x�E�0�ƴ�����^Z��C�!aCmQ�4�a�Y��gF�/�b^��.��-��rշ�X��Y�IFV�N�
ҩy���ڮ(ӫw̞�p�m�{����W�r0n���ٿQ�#�cs����H�9���/���K��N�T��l�!t�֐�����B�]*�����Dv>l��FZg�� �<N��!������%l�~)a�$��۟���&�a��Jdb-
��شU׽�M�v����M"(n܇o_��ר�_�0n�;a�5ݙ���}�h�Q���L}[���=V��˒��=zyQ0��|�(W���u�Yu�<x,���
	���iXM-P���ɠ�s����H*U�!�t:�0��ۛ�{J�p�h˴ $��6P�?J�.��p���0f+d� Ŭ�l�b�������kk���v3�e�N��I����4��`o�|�D����~�z$iX��'��>g�O ��L�����֬��S�q/�ї�ĝw.�����fA�´5��� �����a�@o1vj�\���Eo�bQ��8�g���lc� �.W����������VT�'�w� I����y�����u�1�d��T�G)��rZ5�m�c�����o�GF�A�/D�g�x�g'�a�Hr�����4�g�5U8Ő��w3��x�����c�[�@�*n���N��>7�!�9�� �O,a�T�=&>w�&���2@�a�G��7W�n}�����{~��������${jJ���s=�h[�j�H�_Q��!7<�w���fq,� *������9�Ab��_ME�zlF�Q&^ʴ�&FD=�R>�ʺ�M��x�+�����!i��k%A�$��qл��eEa��+ׄ�j@�t�0���J߰��-?��?ﯕ�@ڞ6�z�祾ad�����z�ľ|i��d,��ż��N���=2В3�Vq3}�=t!x٧U�@�+h����ɷ3Z#1�T�}���w����
i��h�X�L��o�/�`�(A���o�W1�F��6E~?h ��r��Ə����*9��[��
�R�y�Ƭ�ˌT$Y���ff�p�g��&�>p+��~�>F�8�".�6�
�u3�چ�Пh]�/{��;�ю7bE���\����`ȉ�޶*�(C�&�* f��*;���z/\uNM)�R��� ��qD١�!:`�,rFg���6"ڧ*p���J|�\��`��?�����Y.���QX�Tg�a��g�J�����T��*��)�(�@�(�M5��]�Ƣ�����zw��_�)�yd~��U�8�6WwY�.���ل�kE�n��2h��Y�/�Z���43��e%A�c�T��!�`
���������e�伕T�lM��o3���a�H�B�.;�,2w'���%F������6�ݭǈn̦�Ǣ�������,�E}Զ���%{��+1�D��]�C��T�&}v����_��
�W��;�h�������ܮ~ߪ���D���ç��<�k��]�Y���1CB��} ��>�c ��̜������4��G���Ř�7�,{G�C�FС�6��#u���^9�F�B�B�u!0�A�����TW���l�7�X0G�k��E�[_σ��c��������*`B�E�����hj�0�i���E�!��,L��}�#���ޫ�����d�Բ�hXJW#<b|���IwT�ovE�k�Y������*��
;3�!�e�xN;-��{K������t���֨l�0r� �����r9L�7P�s+����&K7��$�NM-~i�#2�OPR����wa�5l��@ߋ'��i���Y��5e.�
N�\�6Uw��\\�����\�m>zr�JU:H����$m5�N|�p�"]lH�%�>L�~��x��U�^��+��@4��+%����YK\o-�}�+�z�R/��t����`�ΑqVs�X�Ǟ��X˨��#���Ik��d]w,��`x��X�Έ��?�ǿ��B;��d_T5,��Bl�:I��k�˫"�~�3��RR�_�!�);�p#t ���V�at��_
΍�ez���NH
����."��h�]Iwx����*�<,�eds�*�׼��F��Ϋ���]f����/�J]�\|���#�#�Mg��,i���ގ��3�`��r��)(iؑ�h����)�ڙ��٪����E�Ĥ7��\e��9���M�:d\G,�As�A���X���b�"��$��p��9�Y��9��2�:��T ���_"�k����^���� ���B�>G$9x�l�9Ń�2(�j�Y!�esb�(p��h�q�r�~
VK]gT��u������1XL����= �Ro��'ВE��rP��ހ��X9p���6�V_%y���z��Yso��4��`����G�"����,���N
<QId�f�gS�civ|rI�BCI~�Ru�Q*���qHM�!S�s�?yL��F�_ri'ߴ���s�Uai����M�c����7wr��C�r���]��#�#�͈�w��u���>VH�'A}�r�F)F��%�@��O��:���+�N<u�~�����K�#�@�*m¨��s�ʨ;TaTxr`�٤�5�Wi����`���J��b��W��E�q���X��ڈ���*ԇ�K$�u("�g�7��'R�'+,�dJ��E~�{�ư$�B<������W���g�)��a��{�'M����9�vca���B��J�W��x]@�N*� ���F�6*i'�t%�XDP*:�ec�И~�P��0����}|����2���\</��qC�)Z�baA�!������*�g�kTJAa��l�HQ5s�W��t��Y�̆遷gH���]��b��0A�a2h�j�*A���'y���S��4�P*%����;�K�9���~�?��;�a�;�,aiD*���-��ãs!��Y6_aN�k�}���_i�B��e����_���|��s�*AEO|���J����c�,�I@�	)��fۄ}�)���О[�����.���SD�M�	=�h\�_�m�A	�Q��e^=�5�55�V��W��Hq�L���g�g��>_��6o��n�w�۱����hfL�O�x����]�����鍚�w�X+�C3�(]�=��X����q�2��4��������^�-�ζ����ܘdrM%�J�'z�p��������Z] [PزM����[��I��^�:�K(手aq��!M�Y����^G�"x��{�/\���[�յG0ˏ|��<�J�=�J6�-� �No�Erb%z��C����]���`����������hB_��q���Yѫm�Kx�<|pZ;��R1G���R����]2ި��-1x�N�AW��i����5���v�����}�'A�(����4z����h!���F�`w���Pɝj��E6Ny�?5\��"��R��ѡq�	h`��y��\I�_`�́=�ŝ)[�P#�G����Gh�ZB��2��Y^^h�%�J4��zn���c�Å#����&2i���9֛7��[�f�&yp��,�x|�0�L^K���#���s�!�b��]�A ػخ��А��<�)�����b�p����ùYp����+Xp6',R���x9+��𙑬bl��j1�ʷ
����I[x����iwV���9��Ν1��m�����dTA�V��z����DD<�ܴ����oJ�����~�g�^wf0~8|�<OȂ��d�_�v�G��lt�x4�d�	p4�>qЉ,��Sd<<5~��kD�Y����Iv�vٴ�h9;��GC`ͽ� �\ng�ĸ߄�b�Dj�T�y �:�B���G��C�;��Ϯo8�`U�d�*���(�[�j�<�"E�`cT^�1x�gS]�AxEN3`��r��8�ב�*B�k��U�	Kk��;�ovҒsHq;s{&2i�*_��~��_§U������ʃŁ��!:6�f��ł�&�-�70j}ϴ����WA��=H^���GvR����i�0�Hc�����UB4}U�ʲN���t��0��� �4y%��AC�AR�!�>���9�樦;Vr��˾t�z��i'	) �@�>�K�H�u?�kPhP�Ҧ�s8/�A=�\V��0[|މ\��9����w^s%���)a�4�W�sɚ�US�L�D�N��J�g� ϵ�n>�/=�R q�Xt5/��J�2�v,�ʉ���؁<ҫ%���-K��(^�M�=��}�<���Zg��k����uF
��ƍ���L���7�w�gvg���x���RN�J ���ɠ��-B����.����Ps�џ�������_3TU��- �R	V�ԟ+tC*:�}�%$��K��]��|��f9G�0�DA���U?���#ӣN��������,�Flo��/Y��	3Z'�\|/����Z�VW{�'���ITA�v#��M�3���Ve�4C�R�sI�1Ѿ��3����s_xP��ӌn*^�b?�l4p����҇!����`Z�ǯJAjT������Qӂ�#7܋r��'I������v]�.�!���gʡ;P;婆���ʟD��!;.`�T��X��m�#.+FW\���ҟ�\]��GPy������w%-����}���k�ݢh�C
H:��Af�+ ,E�u�r�u�: �?�b�Y��M~��}�`Dzf�QF�@Է,�i��n6'�>�˳�z�"y"�1��I��}�r/���cRZB�k("�m}8�5�!:CS.�[��>Uǩ<͑d��.!��C
�-R/-��{�����9�����ŕ�>ei��.$cIh14����#�CjR��FE|����{dͭ�论frU��Z%���8t��ޣ��yt,f��?���ɻ���+d]u	ȳܒ�d�KQ�pB:���,d��������T�<����L�g��`'�����[(���"�t�ļ���6��2��.�*=(�8�%���	3e��H+|��$�;iD5������}���^����8X��^af��C�[�D&�m
�b�P,���Z돼Y�x0w��#W�J"�\/'3Gc.�����4[�6m-
"�W�a���"�CE�����{:ȭ��۴��p�1$]�ø6�;���9��7F�rl@	��Ȣ:%�o
���Je鯗�u�=�.$v��ЄN�u�g����F�������<��^շO��jT,�d$*�2�n�(��I����S���q��i�7)����{'-��>�~�KP
��Ť�ꔊ�ʉ�*�����v��,����V�[������w�VY�����@�5|��4>�vg��n���+D��x�i�K�)1�=�}W([6���$nT��^~Q{�U�K�b�L���:+�ᆐ��1����7�ZD|B����v��(�˭��{���i���d*J�m��c�W��Zg�+�~�h��ߡ+�o�ڏWO�����P7���rall��5�q�J��ѡ \P�bp@4&j�I#���%�?�Rk��T���2�J���wz�ظ_�ww$M��'�Mjص�˟mG6
2͵�^߀ʪ$�Z$��3���CZڛ����~�m\�}�x���?���ѡs`��� _0��l�+�O��	XL[�׭y['�F-w���4e&��4�"YB�V���f�E�o�^��E�*5����6������n�ڑ�ʸ�Q�݂���q��!�S��w<���N�Ǘ3��� �+�!��q'0QU�,I�"l6�#�DVk\�]-ҊIP�D e#�ۮ?�qzi�#u^c)�+ް=u�\��=j�sT�>�Z��؁jt�]�P��l�����H'1��^U�T qj��2��ו���{$���z+�.Ǖ¤>hd�-b�x!D��E=�O�\���]��r1�l�����U��j�I��yw��a8���"v�衎����۸X�Z��	K� s�Ϫ�Y�(���X��?�(�"*Kn��-��%������&��8j۳��)*%���]�\��6�r�^�պW��>IwLBդt�&�r#��;�����2g��t��1~&I��������'4D�nM��;!�;̝�ky\�^`�3q�O���<ϰ;�cJp�/��,J�Z�w�2ǅu�B�IJ��YNg�se� �.p�(�N����+�U�ooU<�f��XDյY��9N��@<�*l9CӖ�06	�)Hr���.[6	�h\4%���ϭ�*8h������ϼV4cT�	��F�ni�|���*��;ƛ�Li�+I��tj�n�}㎌���n.Ͽ�^�R�w=c܉'o�����-~�cLӈ��<D����
�]��4��p?�ؖ����/*l�� �Ia���֕� Q��0�C^�<�.�y��ᩆN�F�o%��G�����d�r~�_c�שx�n��!ycYw�,5?��ګ�(�)Rr��t�H�4�H9:'��#s���ln����nxX_��GG�FLV�K�lVDE%�:ay
Qy�}�`L\�f�
�"G$fv4F{�Q���:>�*���m�+nWÙ���V�{��9�N|S�8=נ�Pv���̨���zlg��b���zj6�hF ��N�vA�Əc�W��A�6U4L]�a�B��� ���V�ZB㘍rT����<V�3cL�*~@��4䏢e|���D�#<o5�%A���^V�dv�9=�;o�%�[,�?U{�U�	{`�\�Y�AG�м���v��/���U�`�����!@Q.���F&$J��N[,5������Ntdޅ���_����`�b�q�.�u��i'�ڄ��?��S��ʙ�W�� )eӇ~�Z��r�柪Ȇ�5`&E��&�+U-{َeѠY_/�6�4�O	������lI��%���k>3 Wݰ��1|O���o�:��y�̏�D8�Я����E֟y��P�0O��jGx����V�6k��B��JT��t���*Ś�-�d�y5.a�D��ǕT��"�T�[�~寁���I�v ��(��-]zH�j(�P�Z�Q&��V���@�� ��WԋI|����[z��4�W�$8�m$4�[	[�%�_�ɂi��:��9G���k�ӄ�u����N�D)�[��*|�T�L�1�Rix���8�ke�@$��+���Vg�:1�Dm���72���I���ޟd�gY�Z\�L���)�rX��M/k�l��i�x��s�5�p�.�Ga�0! ��
#H��u��kk�	��bt��G \6$*2��qxE}Ѣ�`���s9�mK�C���V-�]1��y7XaW�wי��ݥ7�&Fϥ��IO��\!�+ GM�H�(�q�>�,W��x�+^�_�:��Lp�Rl��nD�<@���G���y���5�H���.��6z��f��?�)�n�Y�S���gz�RC�2��z$�`����ږGi�%i~,�q���ɸ��j�=����Jp����s�)ٜ鋳���A��n����X�`"t���-	��4���T·�*�Rq�Kn����{�L)wӹy�F v�P��t�㢂̅���7("Ut�=�I;n���Ո���J��D1U��Wgt;�Z-��x�3�TgϿ{�!7_C�.p��1V�ѶJ �2٥��@9��א�ֹ�6hb"^�8a3A���X휻9�ۗ���.Ň��ħ�D��0ED8>�;�QHW9E�P&��~qg@Í8!�;G��֒#�g��<;����Ϊް]�@jY�+u�*D��/���+���LA�:K�d�Ά�&���|x�+�������{4�����"oB(������ɱ��˚.����ы9��с~q���[�՗@��Z�[������v;W��V�OG8�Q��Y;��ă6ت��
��ؿ�i�x+�^۪�k/�-u�Jq��y�8�:��7O2oݯ����.'7Q�χ��v�ͧ[p�:�B�i~o��~&�,�f�v�<�F+M�� m�ˮi}Z�l�<mE�01�����F��˙����e�>�����r�r	���j�v)W��{�p<�
�?zV�ӡY�sEٍ{0�v��QiT�D0�d�PJ����c�ļ�4a3Y���Mb�:`E�ZС�o�KJQv*���c�amƓ/��X:ɐ�p*�5�9���!l�si���f�4�(�%<��|_|F +&��٣��L���<�&�g��.�S uUJ���뽆�u����YE>�ic%K*����.��n��>C�U��Izse��՗�$���G:���YvGx;�h����EK�
4�kyvm"y^�9d�ݣ�Leb4P�$[yu�d�!�X}�qB�e�<e
���Q�t����!^h��P�K������ �_\���L�E��$���)鰮��/�ىh��sR�_���S;Kp]J�'�~,�In���.��Qbd:C����v�B�D��{�m�f�\&Ұe���?�����|�n{7x��~0��d� ?\'�خ�M\M>��A!���O����<�J'�	ى�������~\	�%�$�KA�I� ��gP�t]����E ��H�� �'���1��Y�dS\�w���>35:q\��^E� �Wwb#���P�jx�Q��%׃�=�|�H?��:�	��?��}0Q?Qv�J�Ƴ9*�o�0Pi�Pr�KMHڮp:�DjN�*���}^||�	^qR�O7���V�:�ɞ�#�HEF�m��	(ѡO"m{�6�>����!f��:
��O��W9շt]t����ocMd��یf�L��,�4�fE��є�����WyBI��􅨏��p\`�a��4h=Y@��2ېS���z#'�x��vń=�+�v�m����0��!��vZ��4Pm*�����I���3�@��Bc�� G���Q��%Z�5��c,�vҹ"X�ݕ@}\�7�Ƅ4�B�ަ�!P���N�ԺX��@)X���:	����УRF��9[�Hb�gI��=�&��'Ǹ��֨#?~ϱ^���SP���ǭ4�/��X,ÿ���1��r9Ht�ů���+�MDOZ�.����"�#l\
�a�{/L�+�SҘ�q���M�ǒ޻�p�"l��\�2��:i�����fO��#�����ʑN�鼀�`;�}:#�Ii��� �7X/u�'��'�@�5�7�)/�<�������b��!�.��]�P[��0iv�/{{�ۑ��E�&F�U�� �ƾ�.��Ix�-��&��	_A ��h1��஬s7O��W�O<.Gm�<9�6/�ժ�:B�SS��$��0yU%,��(�3���d���l��Ɩ�'�;��m Љ���dj�4ՉQ_�!��"���s�bGF _��%�ˠ}��M5�5�X�cR�Db���U{�(G���Y�H���s{U�FgW����g��R��V:�w����y߀�}��<�CH����|�q��7x\JA�BKB�����+}�;�����3�Ee�ޙ &C��7T\�ΧD5C��I��C=a�F'���w�KP :�TN׼�/��l����c�X� 9d�B��Z�5����X��Wkko��;��L���tR�r_~Jδ f�Ej�Ԏ�5y����X*�d�]S�5�F�ak��Vr��My�����z(Wj�,��[W0�y̢j(���m�+���l�TG����>� �@/<1K"0�'�r���͟36h��Mİ3M�H#	mO"טCXʈ��ӿ�|
�ߕ��i!^��z80pY�@Hm� Sw���N���#��9�a���^w
@�Z�6f��Qf���� ���Y��1��"��=A�Cm�����@S��Q�%�L]1+���f�@���(0��O!�O��[�(o��f���;���[�l�����3Y?n3Z�5˜)��N�����~�̜��
�?�dY���������ο��l��ڨR��	�UT�Uv��0?k>ī֖{=q!��н֚���v��^c�6�����'f�M�;:�da`�%�b[R�%~	@��rb���^��,h�l<?�|��L"�.��5j��P6�><3,	��.��ޥ1㶃 K$��#D�^�Ze�D�)j�'��P?���-U'�+5#�zA�*�"�\�w�@�,��2�1��acٸ=WMdR�ЭhK"���9((�Oz��=�FeDw9�]�����l��ٰ�>Y��]�ă�XMM7A�j�Dڢ�*E�Kru�y�(�^�vK�p R0�[ۄ4z&�����7��
&���;T��zÜ��rP+�Ast}Ȭ�yyO8�����`��ô�A���_ҕ��C��H��UAU&�T'�d2K�LNd�Fi�E��<;2᭾��<Ck�0��������Ww~&�E=Fd)�{��GG����w�-I��nZ�5��}��G������Z���(� ��S�k +�P|��Z�0#��4�O�:�2�|<�k�旹sR��/S���0G���yB֙J�l�9y'���yY�b�J�nD�^� �ad,eq��u�*�Z��&�!��d�a�p�������e����-2������G8����)�M�y�s��sU����Z�z4�w��['����1��3��d-�i�%�����#�tB��Ʃ�A�<Ŭ��pU{��\{J� �Ůy~oN�#�|��_5>�|��TA����rI)��sOakKdE["7��<�����,�͑)�t
T|u(�'�'��"8pO`�>�8,f�G[Ip���^��5�g�Zmdx#��P�	b���%d��XG�P��U���X�w	���WX� :�N~؃r�j<�盪���U�`���p�
r�N�l*���gg򕤴�ҟt�B<z���aj¹QooF��
<{��>� g�����*5��n*$u�ݿ�^OOj�9��}W?]�%��)`�݈e
���Y�����q��W�(�qs���S���~�(���QV)�&���'V��������ld����3O�}��F�֩j|uW��b�������iQ���1ݶ&�!� ��Ύ`�A���f/����إ#�o�K/�J�)��&:9��H�Zn0.�'�vN��+�d�Hؽ�\V)��ſ��V�M�Xυ��M�g�����Elξ�g2�U�q_v��6)�[��3�棰I�l��V7��Ϲ+Ȍ��=��Q5y�a���k�aˇ������e�}M.��.���~���/3���}q:�Ｅ��7���UZ5)��T)@աzt2�1
�FO�\Q^&��%[��<9�B���J~��	x�oK�nt�=l�'���N>�Ң���gwgvGL�A�F\enX�qjAL�����A�
?����3<���!*���5���V���+^hN�!]���\D�Q[9�*��hDA=)Ef�6��F۩Ӆ����W�`�j�hO�n�-��zS�.��R�\fJ	i����ͤ�7Yv��Ԇ�ӧ��D�A��oyRE/4OO��t�ԯߢ�r)�� ��'�A0���2F�x�.�n���bӛY���3_�]~̞��J\7A ����P*�Iw��]$����.g;-��|i��:�Fe.`&��B�%=?��Ttڿ1,�[�u��Ex#��ov?F��N]�L{�$ܚ���Ũ閎;��Cݦ��J"ӓd�l�ܒ��{R��M�9����_nK��w�[�-����������w	�]���M�����lַ��8���\�]R�𾸊��2�c���H3|0HA;���K��f�V����+��)��y��q�>���l`�%��O�YB'�X��ѳ=U��U�Q
�'��L�����b쟐k���l���i5`� 뉇�t��k���[�b@�ī���rH;Y������o�c��S��i)���D�u���� �U���ΡR����:C2Z�:���i�}8
��`A`�sW��^�
���k:�HSC�fF�td�+�MN]Q�� �;U�,��"`g�u�:/a��v`�!>��`c�-�O�	���[���0��a�c��KeM�Hu��/���	s�E�Z�r>�
1�<��P����tҔw0��E�i#�
榍��2���|y�c/QܽQ���E$r�#X�V�Ұ;M�����2�w��x�s�H0�J�|iEo
����D��
�V�Bƚ��b$:-�WMC����h��o�FN|�``����0$<�-��7r �O��TZT�BaO���y��/ZV��Jv�H�r�Uwb!�2V�&:���3c�W�Y6K�*^�3r¦��	-�qU�K�;�u��k2�	c��7��3w8usb;��kڙ�čXV\�:r��i= �:>��� H�L�]�ҽ���v�(�=�	���=l2�I�N�% ��!M$[m&Z�d�j��������r�$�Asy��ep�L֝N�\����,3=��Xv l�&�6�Y���1]7G>[��ׇ�5
������#4�S��*C��3�蠔���P�AǗn5�ԕ}�8�]Δag�9���:V�Az��QL�,9R\c,��ހ6"#�)#
��^�_�MvX�/�f���A滔)��\��2 �5G %��"*l����xJ�=��y�u�"�	���ݳi���+�?!1q#��=�Twc䍒E� ��WiVB94Y�q�ؼ��h�B=��U4[������S��;��?>�\҈�l��]e��D� `[dk���+�xd\R��Ѯ��TE���I�غe���ޥ��,�� j�؛��c��I/��&5�^Z|'Ƹ �!�ҡor��nq�(��n��l&^$T�[~|��׆�t��P#u|�m�_�p7�$��1������ϔTބ�M]�����3=a[�t���ѩ.2�j�^_���
S9�	�G���X3?U〸���ς:ks$��!��;��Xے�)"�zYWs|5bXɓ�E�o͙��Y0��0&7��.nb3]��J]l�\g+|잤[G���#U���^@����zPXA��
�L�e����� )����n��Z���{T!C=,ѸEW��
�)G�<�j꫱o�7���X�k��B�K^�?�$�?��)�"0�׷J��Yu~�.K:G��99v�]n7\��#]F:},V�~�"c(kKK/rz�ꤋ��:�4p���LM�<��z;觹�w`Q�J1��ʒ�� *k�C���G ���z����+x�oMX�|�Rn���r�*rG\��o*���T��$�v�xh��xEu�!���7s�jy�����en�R��O^`B-�6�]g;��^���ۚ�Ah�P���'2D��y|�Q;��I!����S8��5����%>�z]�5�8ޠQA�P����Ģ�?��>�T%�v��B沺I����m����v���$�=[�~�:� ��m'Z�"�1tb�⾝1�;�e<Ƣka�B W���q�K��kA�����:�C
�XDl��+Yܓ}�oL���?��I�#H���;9\�����UH�5ǙAoR9���N��3�e�Z:'[�B;Ob�������1�Ƞ;�ٹ��D|�_ߋ'2^�x�Mi��E���[o�ą�Ø�1��e�f(uۈ�Ἁ�Cџ�dnD�(������o�!F��T<�zJ��9�a?�J�U?�5��Y���˷�����HWqs���۳���-V����w��}�1�p2H��r��Nx�ή�d�׃���yR��%�l�����_]/��-�>��m�߿
{: ��l��T"���Yg>�ǣ�=����j�z���+l#����|Y���wN�쮤�<�5T$O������͹�=�),k�5�|�.����HH���?���i,��B����у�U`����������	 ��Q>g1�F���ӋS8c�v�A�'�˚���onr��.ǞT�b�)d:}��T��ظQe%�F�����c�4(��Is/-]&�� :��A���t7d�1���1{��K�q��&��8�xJ���{�F\��Pus��o�㎘��Hyjw|��֖�u��=�s��M�M�s��ź�[~�\���@�Uv�_�X B׭G��-L��'�<O����v�?�(h3̩������I3�K*z�T�_���H����F����`�p2�i�����]��ΐ0��|{
n���g�
</ѝ=��u҇Sg�����'\��`�SZy�*O��5����l��}a�Re�3�0�=*�P�Z�J o$h�������dhN��/�3���y�.$y�B��o|��`޸�z�w#T���SG�	wmӕʃ������|�R�o��I#�Z�4��r�m/?	����S

���x0�4��e\׌ng�+�0�ױ����;؆1�(&����?�F�`��0��ї�+�m��V�u���gġ�#�
 [�nA���F��h�"���-�qw0Գ(��xi��ꚟ}���ߔ�o� ��z�zU����S:{����VNMN�|�U��ۇ��!\쫑�O���1Jj���B����L'�1��HB����`�;
�s���$C��=Mr���9w�ft,�L:����>L�Θm�1��;�.�F�(�G�,ݮ�r�|���6tae��V��d��u�Hfw"ˍV�\��]A(�$�S���yЩTz��"��wٲ���5�]TYD�;������<|�w� ������=��K� ��{��:���?��&i.�;áx��l��G���#"�a�s3*w�p_i���,�P��=�m�x�ȓ��Fk�|1E��L��^Y��޵��4 �M�"��㆓8���c�;�K�eѬ�$�$XHAۏ
����Dh�I\�-�y$�p�E�׍��l�#����F��fR7���FA^�p_x>.����n:���ȑ�����9+��,�c��:��AǄV�,?�'�o��kզ�X�N���+�#Q _�\�d�.�>(^ҥ�jv� �q���x���Ĳ�
���D��U(�x~�n �]�@� |�625�Ml�y#��AV�E�hp���L�{!�X�|�v�D�/��U�Kǒye��Io��et����D������zG��3#�#�?�(gVnav�b��4Q�y��OZ~_"�>�)��h��������m*k���[�>�m�!�	� _��o��b�'���Fn˔���~yw�A��<���.��VO��xW;����x��d6ͦ�Ϫ~��(, QX��eڬ\�P�:> V�2L�m����;h�W�}	�Ï�_�l�ϒ�U�u�,�O?Fy��EC|	8�bE�gY��vaFH�I�
'�{�5���(s�A���櫍}�c�B���Ӄ:ރ�&�m��(ky�����J2݌M����B��[���W����!�9��3�E��RH�"!L�E��[��ܨ#��]���vk�����T�ťy9�#ъU���)�#M���K��M�ǘ}-F�n�
>�i���ޮ\��T�n:~t:9+qq5�^1�������x�ۤ�B�C��੺<r��<����8cY��x{ْٲ�l�!�{Ֆ7���ëƠ��Lc���\i$�j�V\G�"ׁS���d[(�x�,8ŕ!	%���i�ic*�V*ؿ
�.@�2j �m^	tŞ�`��!8߼"t�	�D�n��̝%/u=T����T�ԟ�]��t�-vM9+�)�U(�����Ѻ(�<V��&ح�D���/z�\vB������1y�Wh�C��Z+⭝E���\wx�k��(*=�lCL�*ى�2��d|*�+�cݬX��YQ���[O�3}��O�F/�ɜ��󑽳�u�J�v�k�OCD��7UY�� �/����F��s��ʑ�g9�G[�g�nP��K�,#�� �};�+Cv�la k:xr����i��)�n�F�FeUr{�UJ�)6��T=�'P����YK�N*�V|{$K�vܐ��9pN���8|r�"3K�zN���65�D
*�8�=� �^WpO�Cr���r�Қz�	���Uz���w�t����/>������3�����;��-v�����z��I�d�pp�kjF�����9(\
Ohy�e�Mui(��,,[��1r�g�XP�x��Lh��ڑ�>������,��e?c˲;pe3W��6�`���.#@��í���<ߩ���i�	�6<xJ���s;cy�A,�Cq�A�5����e@��V���e[�'�B�����j�O^%�d��_t�C���]����X��"�><��j��M�%�A��B��)�tp����K�����Pq���17R�`Z,L?���ᙌ�7���ɶ~zv{���
�n�X�?�k̥T9���3����.dY���y�3�V1�1�܍��� J��Ūh],A�O�6, �6nn��'�+ �;��M'C��������u&��z+��'�W�ļ�~�WTbM>�2���
�nX#� r'�,�G����(eF���֎��T�^��u[�|��D�.�&��>o���=��b���T�Mm�﷘��)W��,��>G���G@�[t�r�T���3q���'5KYI�p��=<�[�b�8r�����2�OQX�wM��e��JʙR[S��kk�y�@�T��,��ʜ״k}$B��g�\���͙W#9�D�_n�"ξW&��g�r*Yn+�}{��R�;���J��V �hQ������ZŕV�R}�� ߷�9��T%�����m;� 	�Jy���%�%W�RwW�#��V$fxI�L�|�'f.�]��+�����:~��=*��s�H�ݜ��;���W���)�F�ɳGA u���hI$ja.O�rB�UN���R�ދ�t��i�u���֍pE�hY&�N�P2F�^�~����w'��+ϡ�V��V��3�[������`��M\86$1�Qr\�3��Ly��oX�z�i!Ԁgzi��U7�#�B�'����um��_�1.K2_��$�����2q�����-��?�s�&��D
=�4�	�����W��ٰ QޔcwU��~���Jkhr�:���T��u��^i�|b��,A0��LW�-���L3
��-��Κ��4�V�Y���V.K^�=��zi�n��N��AAaDQ�>C�K᧣�HC� c�!F��G�Y�=U����-������O�2�҇Eq�l��PG�h(,g� $ko�N�a�j�݋@�+�A�/6��^�R}6�>�T�aNX��*eX����CO_J��+q��>�OG�.�e�:���{(
�����\ƙ���	��fP����9	ϔ�����|3b`�7`�a���B5��	ȼD��9�d���X&�u~����C`7��2��B��֣;e?��d�]1. p	��Pp�n�{��-�,�<����"�;x��(���B��/���9�/:�x�8W��@�yH(���SK�����K#p&�� �Ԣ���9�(p�;S`��]!e�{�ȯ%��s7�	�!뒱�/3D������#jN�6Z*��G�^�|CjY��Vn"H���
���\R���^���)��g�}�R�f�y�EXt�;�K������1Ps���]��W�2jQG��#^F���A|Ꙍ�������)����_��ޖ5��~T _��F
��t��46�$hyj�������C�C�@��EQ��7Z�Aa�!��0 HrB�~<G@�o��S:��&���!"���*}
��~���S���l���,�6$��ڵq�T�j4��l~��n`�)��d���vi.kbw�v�fy�0�5�fwiz 1�g�:�Ռ�U��\U�9Ԭ&�Na��D0>��BO&B�0�[��p���]�X�񿴦c>QC�\����\hqx�����q�����?��(���l���0e������.;c�) �q		E�@��|����Y�����rN"b$4�Fe�7(��K��}9���Ȳ���U��I�<쨳�(T��.�1P��4�AW�dÑ�D㢣E����7 Xu�v�+ԯ�W`��/&�}�s�_��C3ޠ�(����|��Hڲ��Z���D�9d9�j �C��E\"뽈�ԡ�"�����!��hڇ}&����ݐY�y�F�݁'�����r�c\�=��������K�=���kFpb>� 61bS���O�"[�	�*�rD3�/C��P�3;�Qi�L�HP|'��UD��6
s��_�[��F�R�F��K�iP�4DM�P&��	�pe���t�u[��i'Ƿ/-i�|qt��^Y�8;�JX�<���F"A<�B��~%w���IUkb�L�P`����ob:���U��H(��M�A��o��=����~�8��Jf{7cA|h��� k���~���o5��Z��`�5�2IH��
!�i��we'�hS�{y9�aLD����h�ǁ��Ax���9d������k��=|�_,�@��B��)���Ϧi��7�5�L�B�� ��l��Z#e�����^�=5�����PR� "r�T}`�a�0$mL���<�M	8�]8�o<�!��n*"���Z�,���
�f�?����5H�̤!/��h��IJMu��������_g?W"0:y%�Q0"�>����ķ#�K-˪ "�Հ�H�-w�0��[Y�_(nL�]$�et#�l�Tb������ ��7䝌~��-+xi� �����5�B�Bv��q�)��,�����c��+F�5�xnp���#l��f�Q�a�៌����o5���Z\���[�Ur�1JSsC�|��^f�
�α1ѫg���N�#��
�e%77�usS|�0��eR�ߕ�;��k"��kg��zbE* $L;U71��#��3����T���\q��-��J��9�*�cw����`.h]�o��q�O�s ��5����KY����J���[�z��xȡ�̸��~��&�"s�WšRv/?
���]XM��!�x��ߗ�*���i�cO�
��$����tg�f����1�a9��z�ש�'�<�;{e��d������d��.�=���������h!=�|���k�T��m��Yx3��`�(���.j�m'��^�u$�6Ȃ<�L�d����
�z�.�_o6��(�
ᑤ��?��y>���B	��>B>��F�9=bG���c�_���vJ;^:�� NG��(��>u�:A���$a�8
1�R��b����7DVj��;x\Q@�*�} r�Xц�w��]����!Ϋ�
��(�3�P����q�wkqKޕ��1������[Ҟ��X�f�6�eW����M�]5�H�:���"Z�81c'@��b��������mt02~�P����aܮ��íV�z[z��*�/ \�*�t�e�ф����V��"�cnm��r�`� ��i�lWO�y�<ѶL��a���茦���㴔t]�s"�u��.�c��UyK�Q�{O�������p��I�t{;����˲E�
��O�$Љ=:A{yg֧���ŕGJ�|TX�����s�:r���ͪb��U��f��+�_H*��3ϯ��1L�Ѱf��{�s�G�*.��P�����ft�S�C���M@z~S�Ժ0�����bX�S�����0)��N`q.YX���)Jv��2��H����i'� 5�h~d�j���g��|#\������=&����2�Y�����G�3`��u�ǵ���((qv�Q$�� �?��=-��D�>|�K�ruk��z����¯Q\z=�1����\�3�����V]��ZXA��0�cc�![��Bh2V&܍ż@O?mm,2���]I�a8���'N#�3��,4�o�fpLE�5�f�y�,Q,�FE�i|
G��� �l;�爐�8�N������5B��:�оwMp~�� ��N;@�:�� 7�O9,�X�A�������)*�'�����;u�B��J�w�v��u�MVIw���f#��vh���
��=��E{���'e��#YHً�Z�2�![)�R��.�=��l?8��L
ӭS���Q�2��+�5���7�$����k)�b�(�1�<$mB���3�N�۴'���_�r���A 5�9�4��?E��+@��VJ|LA�SAt<�k���U��Tz(�1��RB[Ǻܳ�*LSX#�SeS�{5��Cd��h3W��W��O##����|�VX5r�5l���	�����Τ>>v��=��7F��Tj�*?���*aU��՘e,W䵊k��0����;���'�	&��#������}tr8�UƎ*[]܎���O^v��R�x����q��,(C?������1	����J]���I�G9�ϯOK�a!c�M�Ib�-('��|��J���l��d�8K~�B������M��Hx}FC� �np4�GT�0�f�'�7�*eXƘd^'�x���  �^��Q"Gr|�:�7gSu=xk�yuO�/mw#����}��pO8e[̮��7��nlL'�]�#摺���e�}��R,x2�����
 ���oe��<�/�O��1"����Gg\���ZPK����쪅���3�o�p�У$�-�HȚ��t���d�GG-o�EXO�t��� �:�*����o�	��� ����7WH�ޗ��'y����,�sO��A���IAeł6u�
75���G�?�Ǉ�E��0.����K��Ϭ�?<�Q�4<�rZcVr�^ښ8�F�w�6��FJ���ŅA9�CO��j�L��q�{j�����F�n�4��[�J��l)+��q2Z���Kl�3����̒MT�y�u���t�Ƒ�u��]� ��M9m���3��o���[w04S�~��)]����EMC����������n�\Pn?'b����	��h o������-��J�ٸ^6�{J"|��xf�������	P3n�h�.E���Eə����ߌ#K�HɿЖg��j���.ʞ/E��J���c1� #���Ԟsn��|�]%��+��(�}�t7��=�l�ep����ݍ�Fx�pS��3�|K0{��;�q�2����'V�TA`0����ɏ/�*`�co+���.����}�шEZl./C>��p�=�5V���֖2a�]bK��̔��E�a�E���+��>c;��fJ�ٿ�:���OH���'�3Fsà\]�-B�qY�)�Iy�`~�"D�M18���w���
q��zS뻂�"� �<�	�����_�.b���>M��k\&��Z�L0�=�F�aI�� �5�ϐ�1�"���,�~��0b/��H�����]Pd�r���6僬�hw�"~�:~@�3���$�Vj�r��v�"����>l4ãP
ޅC~� �%����aM�6��Ѵ�+0,ܝ��a���@�5�N|ЂS�3[u����)S���]ȌZ�&��`���ZR{�vt����'2Шfo���u�����U��@�h��Ϫ�ډb����1 Y'��n���b�l�2�<�フ)s�����Tl�4�Ir\ާ5##C��
�c�9Vd�/�IpT\d������Q���VO�-[��wႫ�;����O����>��i(�~�Q�)�ץ�#��?G��Xi���T��
iD[�Mh�y�EA�ŋ��j{���J���m�W(E�Պ��&��7����]c�W�مI�(8ӏ��,߲W�M�nƇ����l��!��aUրx����¼�-�̣[ܕ{�HE��J�LdK��r��N�Ҕ��H�⌆�Ja�^����>p��r&��,h�3�o~�k�6�?)�N��H@H�H�hv&�; 7�y���S��]�cY�q�Ml�v�2F3��!�7Z��x��{%0_7�&w�fQ&v��3��W=����9�*f�6q�4w�g]��X%_�{�Hr��q�g(Aa{y3�x��V��;�p�#�|��ϰ��S��2��k�G|c�(�"��|*�bX�{�H3{��c������`:0�f.�.13��C=��FF��p)'��Y1<�S:�^5���t�%qd�q%�N��&�Or���OEN���!!/�x���$_P�fz�u�{�����b ��	��@�^�,~R�>2�[���[�r��ߠ���po�,)�� �s#�aB����a"��m� ��;�����D�%��d
fX���=���X&������������RI�DϿڀ(��q��ˆ�H�I�W�\���(����Y�x-��,����
^+7"�~.�o�JAϡf�>qT��X�Wy��A%hޠ��'-����H�i&���D=@Ny���a�=�5)I�	�G��<�s6��*�d����es�h��ӿ�����`�l�b�����0�p9�gk�<� �2��?:�3��-dPQ_yn�HPF2���$w���:����6�W�k��`3�B�Z e��ts�9�N�'oLCy����|�>��pb=E��PiT
L��h��	�E��$T!2CL�%�A���B�h_��c�ΐ�^[�����?h�RW�v?�(��`��E$v$n#�9�iw@lt�i�S�P��D*5h!���$�~��Ww�()�I��ٱ��nG�
�6�gd�5��~�_���.���N`�� �9���#CNT҅�(��;���D�Y6F�a�Ћ�1[�'�h����J�]��_7���.^�1���\|E=��1Ψtnt]"�m���� �)Jo(�-���ojn�"}O	h[�KN63���\�b�\�0/�#�S�S�Q�$A2\R^�ɉ�^ܵT�H���Q�ɌK5�>� H����ka��!T����t�<L��5Ȧ�ݦ8��_�W*�H[�!�� �r<"���c���bJE��%Դ�Qw�i��]���K|�D�0uƖ��er`����z�y��tE3�~�Ig�pő�7�1}U�����}�QP?�œ���K3 ,g��{o�
{�S^B�#�#�׍�!(�G�R����a|P�}�5Z��4�m[[��vqI��Q�b#�kڼ��,�g�ȝ�4/��,i��[2�9�9�2|~q�z lÇӷ�Jf�Q�>�fG%����\��ѼI��Z��V$�L�K����x>�8*_c�t�+�g|��U/W�9j�h�|h�l#^,�P�f���D����Es�����y��y/(m���¥J�P�$NSU/�Np�����D�˦�}�������`!�7�Z��֎0��`�������m�v�(8�:��^�~"�^�,�E���6�ʁڕ�{��8���q��&F�����sb�S���c#�F�)�:��'�y�������&��b��R�����\\������Q���Bg���X���dFdK}4���&7�0,��>�.u����S>4���T�9��\��v�Jp���7?:#����i�a���U�W��W'�ku�^k�$�<�#ؕ�G-CG���	"H��c���j�&|/��V*JG��C/�.3�%+R<�;j���r]An��M�"s�H+����|�4���ƅTfμ�aj��b�Ӗ	}ymd}�Ҳ$b�GF�+4��εcr�fa�����#):���=Zh��l��b�%���g�B%���?����p���˿!,��N@�:c"x7�d��� 4�
46�&���Nr�ƫH$Q��lj0!,���:3����^z��.q4�r&�u�����-G��m��:P��T�>t�M�rc�@8���0��2��Qe�/obt[�f�[&
��X���e�ĸ-���T@�l�҅I�9.� (m��)5��8�P'���z�~_�7��m/� kk�l�8�����r�a�� U��ò����D�N�|��Z�!���(��'�y�Gvl*W��W���)-��ZP�� ��+�'�#s��n��ʕ	�����5 �Ev��+ii��B��z�#��![g,��#D��휔]�? T�0��?�j�[�~G�K�l�������-��x��T��~ ��`r�)1�y����{9CC�6ů��O��� T�l�E�6�%�<�ћ�7�M��h;	�<�`U/��\�~��ǋ���WA�e����(�*�x�{V�ߴ�"�96�3rJPܣm�f��?�"4����l
�u�B�
�YQ�
8t���'����V�rJa'XP{���P���9����E���c�5MkSZ	8�3����Q�n=QR���q�1��F��<� ���my@�+�f6��l)�>�)���?�$��V��������;jV���kڋ��Z&��/;;�4�&ćI��#Y��!ԒW�0�26]��(�>���s�{�?�H������bY:��/�Nv��1�=O$����xq��A�Y�\`v��s�o5Fy�~�7��Z)C���~('k)��uXsߪ��࢐`"�U�$rueZBlܒʸyٺ�Ľ'温W�O!#��Md�^2�DLWJ�"jD�XkL��7#�ć�����ix���T(��)�g�,=��K
����u\Aa=���#��F�T��Ӵ��i�2����yHŵ��@W໓_�LD�s�:F 4��}p	;��=!$����z��|�q����0��#r2�jQ���@�l����� Ɖ�n��|���R?��7O�
��t)
y֘�a�B;���ٗ��".�0�Xw#Ϟi��%�;���pS�M\M����
��z)X��|� ׯ$��z�x���ʷ��C�:��z��xWv�J�E�uf3�m�rm�Q"��ya�"�+E�j1�Ӭ��"7��B%�|���o��X<g�)Q쓬'N=����!M�7�mj*�B #��=i�����?%��+A�p�XOF�<��MX�œ��U`��H������UO�<��b*n��ݩ������g����<�Ckx�'\�䁉�RhӴ_
0pt��)��\�a�$���f�$����E e.����/���e���b�:�l�C�vy2���� !4��H�If� kR&ۥ�sU��1�FZ�VŅ�fO<?I+;D��'�B�V����;���<�R�8�9mGP`)���G�#�,�&�f�Dh/�y���	q�9��'p�r �I"$xT�9�wɥ������q@�f�J���?S�uF�e{��a�VSt�iM�y��D���W��R���U*����=5e���"��:h�[�� p�r�[N�r�f�+��S�S �:y^�2����V�$�)��Ɛ�?U�6!0Uh��Ws��O!Dۋ�K��c�I��b~7���B���0C0�`��JM���-6���l�A��5k���I�vM����ة��ODy¦w��,6_��ҙ��ըHYؖ}=/oB����؏���^?5�1S��vt�ƺS���,�a.4�c0�zݾۛ܄ � X�dR�CN�}S}O^m3*�=�����s��T�vשC�F����_�6o�t���#�|,���G~����[�?Mۆ"0v���$�m�I�w�c�k�H�I�`|+^���gF㠋er-�Us���c��Io�?�8�9#��	Ã����� �FD�7|By�k�nf�ٿ��z�u8���d�F�A�aߘD���v���RY��U�A���+�N0�#��C�Q�|2�ϯ��_��3u� a�
z���f�i�mi��Uw%+ �`�2�娼���/����8u�4l7��)c��s���+�X3^s3�;��{N��^'
r-�q�����ޅ�m�~�~ٽj8�9$�T�o�&�6��ʮv�Q�����G�vL��^B��sF����1+�S�E�Z"l�=��qZLG�����V+�_-�ֳEt��X���G�;E��&�������ȣ�WX�'�0?>�_�ZM��a�i�D,v�5C6�δm��q�7�\*ҹ�[�D(����!5 %�Q�&.M���9�]�!����]��d�?�飽t��gc����=�U�����ӱ�D`��mk��z�@�3�z�����	G�EH8a���J��:IKZϹ�r_#5\l�q<�*�`u��j���nD�V��wm�'v�r~��D}����3g��s5��Qp�����bV�!._�V+9����˓�c��7�+t�aXT�����+ں�%��r�������k![fE�y��<��}e]�U0�i|ɫh<u�vq.��h�+	JG��J$ �h޸_I\zέ�����s-�W_Ŵ��}�q����+��u����T��v�GB ��^�OmLC��@X!�>�4�9y�\,�z�*���ГI�� +�r
�=���<�v�x���+qNz~�/F����p�����)��'��׍�� ��r}9���� ǜC >�5���5t�W}�8�Xat��/�����@�r@+U��2���N�;�^]/AR�y���^��V8�a�z�Q4+��a���ѥ|���J�R�D)�����f�,�a�N.��<�"������R:��?��g������Gj7F�!OZ0{�r�Y��%��(�qE��'�%yW��A>�z��B��m��,�ݐ�������o���`W���wU�&�whzt!���tw��ӿ<���#L�L��(�HD���}�����g���#]��25er�/l��,���`<q~~�	K�׼�m�l�WQ
x�i	�����7�ùM���H�
"C���0 :V�h��A�� �|#��g�����L����t G�U�� ��"v)>>�w��5�,Y�!��v���W�y�rgt,Uw֕xa9v�z^R���>l�Z��8cv�
w�:��������Pq�O'႙���L�<I_X���R���yڸ����Z����Z��'�N����
�&D��*����W��)�
�M��v�*�{ӽn�q3O;�2طY=� ��b�//.N?J������N=����a�`σ}bn}"@�=C( .�(Y�ġ5�aA��Y8�bt�`�W;iEz��9�^��ސ}�1��<%�(�H������P��'��O�M���A>l���k��( h�[�z>�Rܢa�K�r�I�:I���m����i�����xnu�r�+v�yu��*tA�^�T#�(5�h�5��c(����ZF�a,�^�A�Y� �~6��b@��q$����BG��\�X�e˒��^���X�ȗdfI_��Fă_�e��g������û��{���n<�$�^4�[O��k�/װ�Q�e��"�Ղk�^ڃ�9��s�!��@��BS�d}}-&Տ����E�_.L�u�ڕ��6��-��ɲ���?9vs+gIх�����A#Κ=����&뷥��~߼}�Z��o�������*�e)5n�8����H�p9c� 7��R}%[���-��`.�-�Q;��6�I�gv�i7��X��އ<39�x���i���ꀆE-�!�����b>����`_>)��,1���X"�:�H�\�Il���l,�0i�Wg�-�70�4O6�ZŘ:�;E4�-�0-v��~p=R�]oW \���ӷ��VG�!�R���@���i`���+����~�%P�A��E$(g�N7Jx�o�K��b�V���朄��5X�t���2j�e+���B	����i��Y��<$�)8��@�|����5��	dm�8���U?{-c�Dg�sxk�1����6��t�URM��D�'�v	H@W�Z�2��J�N�ܫpg��"��XW��S�z
Z>�{�ʤb}V�p��B�ഖ ���j-Ʋ(tf@o��-��$�検B�_6q�t0B*�G3Y��u��{�x��g�^Ĭ�����C��-o�r.B�Cg������ʳ�������v����x�1�ܛ_�ȉ�v�k�y��/�u��*Hc6�5���K�%"(a��b�o�/��إ�������������}�[��z�D�$ʞ^����WO�{9pJs�s���7�1�Ӷ��x�8/������OG�w�M�{�xD
�4{F�՜��E�;���	�Д<�"�MK��S��n�]����-LH�a��I���,"�N��5��`�"��ŵ�r����ω��1�&��p}a����
�r��nX�=�-8�\�Ϧ���h�j�܄ ��'W��\.i|���#��t�xN$�PZ�1��L!����fh���啗C��A� 7ǅN��$���J�~E!�`�Z�H���V��i�X"�É���&�&�]r^5#T>Ae�L���	9�ltRȢ��K���"�uMps��
�Th[�4P /�y��o����_RG�sb��d�|�k���:\�
6I�jq�i�sA�s-����Yyܞ�H�|d�C8 eL�xs��#�~�)�^^.� h�d���g��cE.�voh����A��Ct��뽄IUI��`c�%�w�Ke,�cW�<1�៮��P�?76c�M �u5ڊ:�cAU@��c>�Xo�}`y~2�S�hO�9��˔.	Ӫ���0�Ǿ|64�g��%G�S
�]?f�Q�s��@��8���n�H�i�K�V�v��$6��2��KR3��W�[dE��
dP��u0.�o��0I���i#�,9�|ތ8�҃)�B�������)�~Ƚ�Z!�=˽%�[����~��<�\�~���UTC܇T�ŋ[JK�DҜ���2� j[X
'���,r��n����\d�Îٍ�I2���Pq�Y�a�#(�������TI�/`�p�pԟ�����٤*j��{1p��-����Yv#uK��՛R�ϴ[^�I�j�fۮ0蠑W�y���p�Rg�bXt��f�(���&�OJ���=���%"�ͯEh��-M>����qUօ��1Ĭ_)�\�)ng^? �,h��zъ~lWR㋎���7gA�`2�T�g��Wٚ<g�!������(��[�-�M�PD��y�Ab��}�A����B&`�c�dCez�5S�k�����L/T+���E/�2|�y^�kt��B[' ���v�Z:9
� $>+M����N��WB3��]�=��+�_�f�~�O����b�$���&AB�X�����!`.�^�0l*��/�* ޿ �R�~O�x?����~?���@l���S]N�MM�FOJ�V֑�K�c��1ae�X�����T�,V-���k�[q4H��Ԯ�}��C.­�����w��|�Z:�w?R9{��n����y��+�ȃ�*v� �	���od����}�՗��s�k1z�A�5�8\�ߨ��9��>��H��n:7��ƚ�0��]��?Y�6ͷ�l6�B?���~^��0���":<ss��!�S���A���.���_�K+�7P���9'�{u��x��~�K<7	C�Q�:p��6N�Τ̛�P�(����1��}:4��Z18��uP=��@?Ȩ���`!\i�������y巆�YVi��cA����Z!��ւm��l4��8c- ��Q�_��DFʷ؆�1��yš����)B�9u�F�|�kw��/,�����'�ho�g8�͐e�X_U�#7�w�%r�S��r�v!����TD< ��᧟�{Y6m����6N���?:Q���ð��#-�t��i�A�*�Y�S�@�X1��e��78"d���Wk�'�����!��D4� ب����LG��:���֙0ߑ�L��T���P�Ȳ�E�J���H�� Ԑ�X�Q���QX�9K֣Zc��Q����;���t��۝��b�wt��=� ���;�1�<���
}�(��#�&0��<#��"�i��sm⁒��Ɇ͠�H�A_��;aП7Z���!��L�����h�O����7�~[���5�Ǻg\�.B�2��=�&�g)L!�n�y�RI��5�nt�^�un���=�bR��+z�F�wF#��� �䆱����qB����n�6Y-t�w4�$2�<���d��#6�0� �dS�sK��3�`kXX�"��E��7*m��b6L��O���	�����ɪ;�>70h�}��q*@
�N:�F.�j�\}�*���q��]I�^�?fvN^0{]+�p�!㝜�R������eb���=�QAQ;BL�Ͷb�7>�M�|��Q�2�h��hi��6�H�o'�/�)��0��HcB0C&K��u�5���$�љ2�4!�������x�
�tF䷡b%߶�	��)����^w��6B�p�m$��hZ�� ��@���?V��X�2����Gf�u��작����U�_q E��D�Z��w�ud�2j�V�Y�^R��	cp�y?y�i�N8"�;�II�<�~l䵜���z�3�=g,�-2z�n����	vc�-�ԿѰ��W~���J(F��Ϧ4�[��$����fGbv��i��sGV8z�T�eJ{m	sz܉y2<&�r�f�����k��W+*��w����^��<�f+)7�#�����5���m��Kԯ'k4yySx׭��I@{4`4T�j�V��t�aHq/��2��I��b����� �1���{����24��u�����o�+
����*�����W1�g��\L8�Ʊ���8�P#���NQ�}9��8�(�yx�9Lϊ���pp�u�?.�z�EiS0�2�6h��$f2��w�e�	�c
(���sgx�\��鵘ƧO_z�=��j���د	awF@���$'�~Z�-2�5e?g�Ϣl�T�w���rע� 8�pkBG�@hJ��a�=��c�b�T�aL��`��w��P��26���ԩ��Kԕ��W�m� P�1���ߘlǲ�6����nj�,��uo���vv��z��C�j>f�[���ʛ/��V�˫S��JV-p��������"�ˤ� &4C�G����o�è1�� ��ӫ�&�<�v���uA��D�ec���pM�0/wb2��Q�_��p�'C�p3�t9Z�wBǪ�)���2�:�"����'����#W�Xe�`2Ij��!�À�����9>� �۴�*�
W�n�����ۮ�
�Xq�%'��S��eq�.쉜�Gc�jd)��b�3$æP�`	��u�����k���\��yopqp��(��_o7p�U[M.�6��E��|�*���}e(�k�ԋ9���L�~����!wxm(H�������7�F��J:�r�	p�(R�$/�x�9��:�s�k.΍���-KRj�jFЉsj0⠈Ҳ����c��DB�ܬ"\��o�o�����M�~c�X�\��{lzTŢ,��.��n��O�Af��h��KZ#�6��� w��Ap�$:����5#tԒC���q�]�9s��bNP�.z>��Nʋ�7"):7i��&~��%�rˢ���{G�sv�L�37��W��,�y�)�>�S¬��w����t�K��T�fb�A�Xi}4=B3Rь8��?YE%���zt����E�ڌ�޺�e�*��f�����w�^�♇eV���1���Q6� �P� >b�����`.yb�\6'������ԍ�ғ��zR��u�}v)�\�:5�����S� �Y���v�U8����_K��$x� �nW�3bc�/���ӣ�����E�}W�S%h��j�ku���ր�+j�{������Q�/�a6��h��uXB��c���'�_3ߞ���p���E��G��s"Q����TK]��ʹ���F��}�J�n��$~���F��4e���+!E��K�$w^��sv+�$0�e��(N��ү"\�h�%��V��E��Q��,���ԯű�Ig"�V�W��Ȝ4��5�I��;H.�_{$��s|P�-�շ��@g����q�ʠ�/ Ҷ�R���D�j���G,(Z���)�=֘<�O&�Ї4�8���Ӊ�P����a-���t�(����Y���7v�Mt��&]�}�u7c�7�Kߜ��y������\�Ns�TST�I�F��[���Pk��5/�X��\y �^����m�t���_�R���T[�? �c9�']���|�y�;����FS��QOQ�+��wlM�	��sf`���y�lXӠ��WZ��$u��{�T�ek�L�r\�/酛~�B=d�����1Ps��c��svi8��V1_yM��&s�"��Z��Ay�A@*M��̺�W�j<|X�/'�KK�Ғu[Ui�G�G�)HC�Z:�� �*�J�t���oE��Pߴ��#nށ���$Z���W�F\���R�fD�&REw�H<�wgU�d��F���jFKO|T��5�K�t1R�	_�3쎹Z0���AƩ�ґ��S]h�Zx�A�{��q\�N�0�>Y��ƈh��
���A��!�E�L���������;�
�W�s(N6�> ��*�5���l����mV��Hf�mx�Xp$��J�������N����5
�8^/�>�P�Q����9�&0S�,P
w��p��(M�m�
�<�L��ʂ��������;�!�OV���6��A�-A8�T���5āR���ө�?hWp��.~��5�(�1=��Z}��M7��Ԛ%����}�S�8Ā7���@f{J�{Ǆ����xW� �y���^�Jي�ۮT�n�ڑ��?\5��T���e3R��U���6ᡜi
6
��f���#!�0,h����Ҿ��Z�2H���޵�� 6�d֗���/�w�"v�������^��*ə�"�C�8)OӮkT�uO���N��~����i �\aؖ��w�Sj�x @p��t~�~����KA�?��T�%��F":]� ��?������ך��c�j�|��+QZM�xpu6�򒸬�o��9���w���iA�N(��S���
yp[#E���Feo-Qs܂��?�L_d��c�ֆ��F��:���]�4��Shm��c(t��au�	wr��|�y�APD�M�#�$�Q�T��?I��%���(��n,�!���iS]}��3��<��k/g��T���� d}S	�SvC��f��k
+/Ӎ�q�����Lpܫ��e)�'ީRO��rO(��|^��ɫ>Cfˉ	��Q���8��n��~�X˨fzn�W�������.�,t ʂh\�ƫ_|��n�bz⏆��7��(����Wh	W����2m1x|�u�%j��a����tT��0Ι)Jj�UB �'��@͂�3Ԃ��a��FA�p�� ܄~��n��'m ����,B��ѣ�e�d��9��sR�����8�1Q�O�|{҈��q�7KJ�#b��k�s����^��dʻ���e�b<M�t�3&����o��Km�lA�A1J�ib*s�p�����d �֒�M\��	�y����U)v��"�W?�Q�Y�ϐ/uw�[b����1�(���k�^�gܵ��0oS%.ɷ~	Q�(k�̈洊U7�����_\VqQ�2����i�D��#�H,0Ŗ�m��+r懻dE�,�*�����]:A����|�Z�8�;ט�(��Xb�I_	뚠�2N��.c�N�%sx]/Vn�:.V�|]��O�U�GCUL�i��4+H��!}��F߶#�xBZυ�"r(�[w�i�.$��u��w�)ؤY���Y@�ˬ�
��pl�Pw2��V��s�����x�v�Q �Fh+Ÿ�'r���_ή�a��d���w$�X�~ʄ�}��2NԖ6�|s��u+ >��P�0���|y�0#�2/)Z�l()�s����}����l����k��Y��x�?(B�e�H�g��׾C�S���]��I�Km1�G %@q��J�V肵�X�;B�ۈ�����&�E��v�{=�f@�^�{\v�����.dh�&���W�>�ԝ�?���:�Z�����v>�_I��k�U���9�8�������O�y{҂5������^=�:45�w�b����coۨ8V^&��%e��m��q��y_��!$�Z{�gef�Hz�X��9��zA�������"�+%T�9@儝9On~�|iu��*	�UP�NT��|�0R�i~�L� T��o"��jRsNm�Q��Vk��m�z?�0p7��[��%[�6A9�1bId��e\����~��(~��⩢~ڡ���4f}����xe^��>��pǽ]�2���#?���.3��Q���PD�j�z�uT�='є{�:��͎*-_�Wx,-5GJR��V��ot�Ë\�*6�mЁ�9�Ӹ��+���n��Kmd�@c٭��0�Sд+Kce�΃�g��B�v�����ؓ=��B��,m�Od���SB`�C�ä����|�I��q�I�ճ��+
2��ӄQ��|���l���Q�V���/F�c�y�>r%?��";�_�n%��p�N�$��y�~Je6ݙ���w�����\R�N�c�/_�GxQ/+蒏z�y6t�*j:�w��������uגR+�M�^��Y������:���ψ����f���2���M�p�55�6`xH �������>q��e;�
ؒ�4/��|����o�v�"������O��)�?̘�=	��+�v	�M��D_sL=�E#�E�]�Wzt�F�.ͤ�$������J(����[0c>�<q��kmr>�4٦`�ۢóè�� ������l�P���_s�b��s���b�teN[�|�H��q���d��Q+��������@I�+	�������l�N�N:��.8(�2��U�n�����Ųp�엽������%��W��@�X*��j�YC'[�q8�g��f)��,�iBo��RA��6�u,K	APoЯ�nV>q@��(I�M�#a�؀L�4h!�e�F���E5�H#�f��M�H� m�k�B�T�3�"�P��A� FqÝ,p��y����%#��v�����"^N,1q�Jդq���{"~�Q��a�-0������8Gr��/����:$�^n.Ѧm<�����/��j�c8b��ca=!��w��.�$-G �{�S���1�۝���9�����Qp!�Z&V1�Qt�Я5��N���D{���k�䷟�j�ʄ�83�������o�5��Dud;�f(�>j�@MNbG�Ie�\m�� �1�0.�v�B��
�2��7�?g��}��BF���;����t�d�&|���i�_��V���h�!���^=c��A��e��پ�x='����Ǣ�4:�p�pI8������֜y�o��cUo����1a��61��c]ƿ}
�W��V���bb��%#=Hn�)y��-�����1�AB~,t���m���8c;S��)"m����x:oTNm?��`|�������_����ʾ��mZx=n?Iel��?R����@����n ��&��F ���U��ځ���z%^�c�Y�c���h��&��NΥ!�j�����K������xّS�0��0�K��V�HD!/�/S-�7�<�&"w�c^k���I�P�a���B���>�7p�%����3�ʯ]z��u@ؑ�X��ƭ�$�⍇i&P��[��������j��dz�0�D�/F��oL~����O����L���~��>�x����?�-��Ξ ��r�2j�)�z�T7	)�xv���)O�����B)\a��D��ʕ.<v��&ۅo�cIJ��J��i	
"Ҙ~�#��_x5=F���δ��kS`� ��}}�:��G*��NʎO�*��'��[�8���.�JP�������3���i�lv-��kr��O�YOΜ2�kT�	G@i�r�����nJ5q>���/zI:P��H��A����&��@�~Vq@$l�Ҿ�|��g�y�T���f��A1����uBN�`z��7i���NMx �[�:�w�h�|�NpW���vD��0�J,����pu�?��,��A�p@�̙�w��>���N��W���e�d��X�׳I4YƂ1����k�s��ϢnB~�3�z{��|��*�ĝ��+��6v�7I�f�MYXlV����FJ��ݔ��EI�CrD��b77�'�1�TĹ�u�֞�9���A���Bn�� �v�0$�*��,���Aw3D"����[�N��$7	&Ti�,��3�����_��WV>�D�H������ԙm�"���T͏w7a�Ȝ��tq�����ՎqV�Gŉ� k�zI.c�Ab��Ha-�z��v9{L2�Uʦ$Fa�̕��\��k�Z��_�-6T m{I�W��R`{���H%�f���{P�;rr+�ϒ���֒�s`�+���qD�M��OY�|3A�)쏆1}&�c#�u�
<h�K�R26��W��ՅW��k��'�.p@�:�m40=�ŉ=)�X^4�/O�fMB�D󐚤׹���Euӣ�E��=m���7�GF���k�Iܙ������6e�p�TY���&ă�9�S��S0�gSYE�7{��#:�J�v��W�}�s%��
�jO���k}e�DR��%澅�N�}��]4:K��+�1$u�m�Cd�XĢC8�'�ʛ`�����;�T�~=e�Z���:��wB���[h$M3��͵�2��6��ˈ�%r0y`�/Q����!��f`�q�R� �F�A�����4Er�9�Rn��P<C��?��D]23 �J}�ͱhOx�~�1�e_Z$)[#�<I�y���Y����ĸ%1@�yo=���v��bl�k��j[�I3	_@^�@&�����d�k����U���?���i�r�3P��Z�Ȃ�Ơ���:w�"i]�lN�#9��LϜ���^C3n*g��~=�`��%�o�$��_h���s9����Q�B��jo�0�Q���D�=�l�}	��o�ɰ�0����#9�^~��ȟH��*sL�n�?�+�}�.��J�2�m�c	���G�q�!Y�������\��~�SuQ/	��=Q4�%CiM�����͠�i�ܵ���{�X*~�*��[8��E>�5Q���6��Ad`�h��jȇ�������a�sy��c�20��΅ O�{$���J�o�
�kB�P�g���qIϐ�r�	��-.�f��
tֹ �p?��o��L3����F�$`ɩb� �h;r|>m!��M�1Ԉ?Br���Sy�! ��3���eF!��YF�!��Ƈ�Ļ���Z��dq��E�QJSppP�/��|4��V��+]YQ�i�p9���;ƱpsM� �!)մA��  ��
;wo�a� ����1^`,d	;3I���*2;=O���D�I��6-�+Zc07�[|��U���W��,�ș�k�+�p>�h�!^�i�yƝ)�<��",/ݬ������u$B�-������f,Ļ�N��J����,H�#&�H�X�}oe�Nl��c��%_��L��)��h��^�xoQ��ՈR�+���.댅��˧�>�Â�X�?|P�7����8�[
]QkM�ۖ��T"q�Y��u�S�T�
F�����1�J!�sE��n����R/ʜ|��\�1O��g�����+�{Pq6�𺨀C�ފn����H @t�=І+	���`R��q��&:����^��jQ�Z�ߡ�%z^|1-%���\��V���bl�i���F�j\�c_H@[a�Co$."���8��T������{b�-(p���I#{8�?�׬E�h�#�i�Ƽ%	ԝ{l,�ee"���8�]�g�H�\ENRg�\ʥvsI�$��x-)*U.[��{���h�B��%�C���wB�[=�Vkْ������5SvgI"�sA�r�b����%�i �o�7�S��
���-G3F�wE�07]�&{�p����eѹ�V\�Z���ϲiGo��<TUo�5�\Pj�6�����-o9#�j�o+�pl����;/Im@"z��oZ�uQrW��b��&�����=o�d�!�I��.���2���ϰy��N�S��v�8��8>�m�<����c?K���+�B5	g?���m���{X���Ws�b[ӆ���{$?�^��(&(@��������~�nkm�!�&X���u ��÷��;� 䦵*�#�
��5���;*h�����~���%n��ڡ⍉2��Pc;_�y��fJU�6������4Z'42���Z��}G94��oj4�0O>4!�3��+�7�ݔ����<T�c1.`�-;���^;#���Z(�֤=�1:4�ʀd(����T�Z�:ei���M�t�P�j�x�q��z]d9�m�Qن�606�������4$����uM���;��4��{;��גO�P%��B�$���;�F���c讙Fi�q]�Ut����l��DX$����L�c0��,S�S�`n@�q��Mz�	�>��|)��uc��;/b&�\<3d��o�豣���E�%��W{��ɡ�F�8f�~����u�Jxdj���g
(����[�D�Q�Wym]��Ҋ�g�z*��r`���$���pnb���'��L�"�{9�W��;�u�'�DV--nc�q��U��y%����٤�����IL�
\Vﳑ]d�����e9���3�.�<A0�4s�)!ۜA���jYV��xYr��7�p����{r��\�� ::�ۥaW��ZT��ɉ̎ /'���x�������߹_)GE�;�]�N���89m�c>I)s��:�Ynu�p�_'s~�k��'��^�����/`�\2LY���*1-dW��+���Vc�|ơfMP��1v�']޳:nf%\�" OʓH�o�=�Zg���xV��F!��yO
���ߟ�o%��d���C����R���b̞���/�H�-�
�/=����ED�`
Ύ�R?�����[� �O�A�*�~|R"į ��@ZD4�ڭE·�`d\=�k9ty췸V´��c5,�A�Z�>�Y�<f�[h?<v�3��W�ד�Aċ3��.8��M?������+�TTʌW�0-�PZXם�sRe=�D8!3l(0]xs�__pfg4�,���e�/Î������?�н ���_*M�σ+�����x���XOk�	/U������N�Qȓ������I�� @�C��Y�x=m����)�Y:(��0f��"����_ۇ/�d(�T���ķf����["����z��h訕nt"����ɒ�E�c�a�OH=�w�������T��,�=`%,,��L���T$���&T�>G�UzŗW�Q�8�U�BYi`�͗_�0թ�HZ�#|���L�ù����_,��v�/1۽�\�G��0���)����kg.�iSb{��o��=����ʹ��Lm������ݯ0&�g�5�xw�bk�Y��G�K�g��A����1	�:q�]�ۭwlya�+�l*��|���&BnO�o��7HP��Bd�`��}^� dU�#����oQ �U֨"�6�����%�Q�����I��߼嶫��l�H��%DU����C_�&��Y�(���䗜�����* `�u��#�B��Y-5OF�&�i�G�.�%O0hq�]�窀��y�;C���X6��w�(��?Q������5�7-�~��[��[:���e���7�2^�/������i�����(�v�H���vs������K�Yi_�h ������'�p?�7j^ۭ`sYvq��dn8o��AfDf/gl�zPWҐ*�r�FT��Ъ^.t���� IjrG5+Z"��?X^��
�7+��nA������KQ��ʅ������U�ѩ���}�<T,Z���2�+�ɟ��=���T{%�>v��HI���akɫVD5�࢞e����ܶO�L�o?j�n��A���ޟ���q��\�N��*e�� ql �%,�ˉۀ�أ�u������F!��="�bP
q�x[d�[c�(�D=^%�ϛ���h����#6�;nV�C�a��L]�>K����N>�vK����B�w�.r�<*�L������Ϧp�2���|�I�������x��7�����#�qU[����WZO��+Hw߰v!�X�<h����di0Ƈ 
'C���`�
�-8�l��$o9�!r,#�K`V7���Ac��|���![��LXOb�6�4��A]ĩY�s����T�z6�:O+�%�UA���M��b��d����q��Et���)�'�1is�1�캉�W0��qWb�y8��x��fV���g������vӏ�=��p��Kc�QO��e#��t���r]�,c��m��%�9��)�Ք�D��Yx�hL�ۗ�����ޕfcn��V��:����*u�g�?�
�99������6�Ac�@Ы����o��)F���w�@��5��9����,�/d��Kj������XH�c����$:������a^E��,>/�R��U��i�kXxK� �i|2࿗�TeW�ȓ-��ӌ�f;r����Dw�Ol Y�M :������k�0���=g��	���󟹀x�.���w�m�ͽ�ı1�$L��!�!!���*��l"M��N_{[Q���.=��8��,E�����g�| g�`\�W�j�Go�-��7��/C�G]�dߍ����KN��m/H�H@�#h���k*h>���s�C��;���R�h�,_ ��*1ܬ�rE`�~�����A�S�r��$��#��jǒ5� �&�~l6�K²����_1��6s��OVP>����;�5�2����V5�ui8�[C��#�41���&K�^׮�T���.�IW�v;��|�g�[��ӓ)��V�3 �Mc��PL�W�q��Y{�z��,ݱU_|��O#F���V��ha��`�*���'w��M?_ß1π ��z<�K��(��O+;�2[����E^�#�d`��M��pz����?���f������繡y�3H0(�
=1�Ɗd_p3��~�TQ�K,ƾ���\���!���W��1�E�K9Il��B��mz&�lM�!�~*�l�v��):��9��I�� ����iԢ���bs������Q�+Qu��b�:E��e��\P��.8 �a:)E�iG�t�r��V��J�̱��Bɜi�*��<kb�S]4��Q[ם0o��C���u�j�|P�L�An6~��Ĭ�!�s��]��Xʉ�Smk�{ѹL>(u8��-2�/M��K��2V5�{D7B��"w ��H����XBg�R�h�1�^c!3%�f�9�.�ܐʓwu�s��q��թ�>��ƥ`h/�ѢbU\����7l���p����6�)��;<=�`8���5~F�g5�5X���1۔��D��Th�Ŋ���	���\b����4K�<��P,#���j0jo�o3#'�)���a�2�yN}/��4�&4�G@A����/s���$3�h�I���mOP��9Ń�����$���tB������u�Mۇ��n�9l�#�Y�Wי�Z@���ӽ���U��=l�~�E<SЂ�
0|�d�y0ն�E'� ���\�9u��e�kx�i���$��Oދt�B%�'o������'���u֌V5A��++�\9�kf�_3�_��T`1I���� �Y�e��}$Y9(o!�5@Ŧ��}��O��1���|Hmnc�(awMxKYp�?��w.�b!H�����=m���ƖDW�s��|�<��-�W��o����Q�*�s���>w����Ӻ�儻}ѽ��D�NZ^�\��%��y�l���}��+^�� �q�0�a�^)V�,�>�9�ep���Hl�%����{<?o�Z^L'f:l6��;��t�z���T
�Y���pX���1ݔɷ��G9w+W��g�>!�^0�J[`Ԛ��s��,�\�T�L��Ի��?��r�ɷ���r��4X*��Q<�5nr����5	����>���A���[�j>e"ӹ�h��\{I�l�{�1BTn�]vHn�gD�~"��������e,?��O���lC��Ja�wܹp�V�m���t�����M�(g�����h��)_dN Y��e�
3���F��{�*�c[{�5_�� ��֏Hdw�A`���\(z�ċ@��a3Q:9PYq�79�a�2k��*�8�$�\�)�[R-�.�ƈ��3��m�5]��h�	����e}�<���h0�����L{��$J��x��X�2 �뻁���Q[��!*0���y� fhQ=d9�v
@xn�pp@7��r�����͍�|!�Q`<Po�}I����UF�
M�:-Y����sɋ�<c'��pb��,���$�q�2yrѡZ,�ǞWb)f� ۛ�7ݪrjB�(��#!3p����1�l�&��)����s����U�Sh2�y'[���s�γݙ�v��S��Q��Lړ�i쮽_�t@�<�iyˎv��#�ۼo��x�9����-�Oa��_V�A�`*������}XP�o<l�?e�r���`�в��f ÜO���g3��:]C?�̍r�'((����<!�EN�Z'��2���/��V���r'��v�Xh�J�|�z��"|`�;���'U�xV8>�S�9��A~�Ab�%f���Ky��T�OT�-����K�D�	�q�[0�J��\�F��(u.��%�NK�b;"b�k�F�p*C�Jt�8T�R���W~�܎e�7`�j��b�wqr4��|��,�hi+�]Q-� �ɦ�b>�ײ5~P��S�u�ϫ8wSgv6wj�/	��yy���)����b��:� �~�hW�={v	)�����y�n ����2�qZ1|����WY!����K%�9lR�]����"vyB�W.�%��@���cK
�����?���R}-�$��B��2c#�R��a��:�O\��ˮ�r>��
�'��z�4��+W�ɥ*�0\c:��Y	uh}e�O�h{,�?�	�3�Jglq?U��ba�ee�{��	j}�8Ykߖ�L�H�ޢü�뢒H����a�|��~�!��n�O}�M�!�z��q�� D�)m+��,5�wC�ÙL6]8�ΐ]�«��rE2A�9����n Q{�*���_��N�%t*���4��ff�t�J�N�ꤽ*j���f��q�x~��F�Б�CF��d*�dߍxF��"_�j��qnV������[JW�o���,@ɆK ����:�*-@�(�
��Aq[�	�8A�+P��]0�,���W29���)ٚ���RiY�K\Z�w�zy������=��.��.�ssyv�����X�|���+�2k����X��r4�)��Zϟ�*z���˗m�uۆ�����ɦ��K$u&�X�n���ے˸���)N�hY����hMx\P^e��ǡ� ."��%�͜Ao���4��#�?��Y�7�T�J$"BN�QO_6�]Z�@cw�:vQ���1�c�/U���}�%�M*{H~X뤏S��tʍQ"j/�;`��������je�+�9D<��o ��VË�E櫅kG*#���T7fB-Ξ`4n�o���d:*�6|׳�M����!�X�}���%�P�S�f5�HX7l�0K6�2M�'��YG�]'U
�;z3�ħ��p��Brlby*�O%[�p����]�|ۓ��$t�̓�l��nz��@�?+ f�]P.ǲu�8gT ȓ�x���m���0@���!M}aF�P�
"�0��-��� ����1(��#�U�!ĝ6F��ji�B,�`��k@��~��G�['��m �{n�t{S��K�B���h��w7F��ؔb"j_���%���7�M�adW��f��eWu�1+ʧ�ă A�$'�_���aF�̛,$K��Q#M"�6
�c%<�l��Ջ1��XŒt7�'@�<�t�N�(Rp �N
�&��酏l��$A�ո�<��+�KZ����H�s���	�3q�����6�|_�t�/6M�B�"G�9�_��4&X�c�Y3�á�\����7p�?/�3u\����G�O�td�S�k5w���Q�#�Ϣ����e`N��h���.�2��;�.'�.5�z.�&��xu�l>����Ͼ�z�J��'!ξ��6�u�5�w�A��yL�ƘM:��8^R�51ɏޝ�sE��Ji�c���,�fn�����>o���A��!Wk0�����Nf�YN��޹�[H|ؐCkZ	�εl��߬����c�y\�]:�+�H��z�+�I���t����W�|�D�pY�X�}�>
ò�)�YdB�&���օV�̾���R������.�cGS����P�\뭢+긼�
�F��~#��g��ɔc�Eo�3���X�\8��D)ǒ��xQ��h+Gq�y�@�e��bLR��M�W_�@�㮤 ��dg�h�R��:�+��5mT���ϡ{���G���mc�oTN���õxl�F?LE8�["ƌ��0��أ<��B^���t.X<�`��W}g��Dm�y��Ac0a5�����F�X�D�B�"=q��CYX/efN"SgId'�r`$���7�@�m"1k^sfxh�޼�zD|��l�(�t�	������gC� �k2Pi��C&4�hħ�9�����y�ix���H#й'���{�&X|�b���Wy!�K���K��B�E�4��_��fK����>�"�O3E~�AX#��ßy!�hX�vߤJ�h��hc���"�<ӅA��t���v�bb�������<8��wło���� \�ψƚ��������#���v���U���^v>�O�-e�5���&�f����C�Ăh�:SGwX��\ǜ^�G�$S�l��A�WnZ���G=�Ŋ}=�� O��QWݫ>���PD:)�5r6�	W�;v�!�븊��'���%G�ΈV�U_�O��$�	]��¤��!��;��:(�&�[�e;�y� �F���{���	M-Q]1m�u�l<�	����>�.�Z��5�Z�9 ��T�}���v�i�
�d�j�[��B�2��;�Ro�Д0<��^��8#�^ ���S�g!���	�p"����&37#y����כ��H_N2u��%U�9�9�6����bE��h	;dd����T!�Wt�IM	���E�Rl�ֽ���.��9|/�qq����b��$Z_/��q�����(�nO�~�(2�YrZ�����%:w/�1蘭��ͷ8�>?��2&`H��Jּ���2Ai]-��*dr|����.�~Q��yǗU�QI�����cm̭�ɽ+�� :�/'��hX�S�&t�(�-���V�,��Ѝ�b�A�u�7��~�ȸӜ�6&,S���>�����U����K�y͞��Ë��?�����!��R�Lg�4�L/���~Ϟ2K�s����=9Y��/4H�Y��!���n�Ǜ<<=�7���S?t���W�4����(qk=�Z� �4!P�=9����:�Y�	I���ރ��><~�y��Y��il�j{�E:n5��ѣP>�����<��F��$b�!�	$L����Zc���x��'���RzR
h���7���5�BV@,��+�=��1T���yNxP}��U��V��+x&��nI.��>�=ՀוּT+���#�s��Vx�w.BS��[BW���OxX�r��,qk̪x�[��cIh]��V$0W�'
*�|��p��t�ƙHsz��?�:�f2����Ol�FNL��x�Q��LXY&���R��{����X�s���q���1���Һ0���|�3E@��" 3��y�;���X9��զ_J���L�όO��h5��>�jir�8n�����`����d��U/�����(G��@��JT��r_�*(�l�A���x10�!%�Ic�W*KP��"�\��Sf!���Q=z��Yz&��],��LJǔ�D�)���2�Zͩb8/	�J�vn9��3�Z"����Ek�R�����}C���� XzaTl(�ϾO�7��I^OFk&	��t��rJ�M���x�D�ool'�~���T��·���\v.*1ӻ����A+�;7�l�zsa���#�~������Z@IhXp	?R\��܃k/�xW�PE�͒�9Y����6�=C��,<E�X'�
o�B]-�����Mu�ZMτy���̨r���\M��M.�A�FY0M���N	���s���}&�p�%`Ad��|�+��U�T����/{ݼFEk;U1q2Bj��îܓD�sgU�ᣓ�E_W��p�W���R�Ϗ_˳��0���xsR�t��-G�<���	j�-���$����[�,zGo7�g��)k�1�4m^j��+�9�	����a��i5XR�"x��pF����0�B��iG�>��# d�o/�����H�H�o�!EP����^8��%��F�'4=wQ���0p}N��{V,h@ &�PTz
ܾ-���jL�氾9L�ӂ�g�]�A�ʁ�`}��9�3U?ڂ��g���:���S��5�Q����G@�!SG!�Wܭ��ֱ=��Ƣ�>����Y`Uh���oN��\��b|ؠ�z
j 8��.���Do���O���acq�p��ӄ�r���%$U�����n�ѡ�W�3�w������>1�ke�ͱ��<݆����^��M�� 	w�]�~����B��[c.��ny^�:�[�o��7���&FQ���Vu�|�X���Y�@����Hx�+���m���Riy+��B� fW9�0UEWxYe��!X�.QA7�5!ؐ�.;AZV;+rL1��Z& �_%f�O��g�h��v ��\E�jjG���	{�Ak��q<͐��Lu�������Ƭ�gD\�?s����g��z���0�@��x#??�3%�H���9��njg4��@�4V�n0{Y8�o���lG	��xj�4��-?��z�F<�"ƌ��U�g�����jI|6:����g�X�8槤�c�3vvة�.�!5�O6?�z�z�M>H˝��:��q���2�����`s@��FC�u��&��K[��� H��Ϊ|�dѯ�P���7���1T{��_(�����S[�@��I��^���eң��KQ+H�ꘖ$���S$�C�Pq��&�C_ �rk�%�Tnv�e��Uw�0 ��*�V"(@ O��Q���a�/��F��~�6VK86���#��Ƨ�u��㴰�O[�X>�����9�����e�O2;����2VD���"�OeJ�(�NP��l?���n�ٹ꼵���h��LE�\�X�_��Ye�L�Oq�ܡ�џ�;Oc�M M��Y��N�>\~z�m���1{.�%��!�U�H���	��|�(Y�M��Z=N��(�������>�a���ne�H���3���z�w�ŝu!ÞZ�DҐ������pmK��ub�d�e�#��6U�C�Pxh%�1(��S�����C��#�k�E�q�C2�f���<Y��uKV4�fW�~���B�Lډ3R:m)S���_�-S�[�~
���*4۴�
�B��-��*����3@�~�BO̋_���ӈ$�g�tK��k�O2�H;M���`���D��F}Kr�����XC���R0���_�}��, )���su���/��;xu���o�k&c���4?
f$�`��*���s5����i.z2��!M�%�)���6L�2�K_Β�s+2�����$Q^��`^T޾��*�/ZC�����n-�����wġ}q?4��!���[��'{.���xcĉ�52��L5aT�>\���N��������,LuM��/�`Hł"�G8���G״���$��DK���h���Ku+=�?�* <�gy�WdWXtq�V����wh�0�&ћ��n�8��{��d�to�bas� ��	%�s�理���ϲ�椅o��C���`uu�������nx e0�Cu�SV�u��}�1�f�Ҷ���;�O>�g����A�a�q)3:��V��P��ݟ1��^�(߰.G�dw�,�5q|B�1?�A���Y��fF�EsI��C'7Jj@�j�8�\
[��l�ͽ��|��>�n���B�x�"��.���	=��qk��dR��?��WaA��ذ{Ԛ�Ե�m1�dKw�S�����)=+�^|�\��J\@-�,Õ�J��;)nG�*Z3J�����"aIEqJ'��u���/�ꊅ\* >�i	��
���P�v���]��#��:��H��$�!�8m"!�jx#��1֢s���(�)7���/R���F|4�v�g@3��~,a�T&�ҹYVӐ���[N�Bw�jQB�g0�!x���f�d���?�Ş�/h����t唉�1C6
 ���O���E��B%�9�,��� d��������c�c�mP9��Źa�ݸX�	Ԡ�>(ɱ{�"e�ơ'��w�Ԙ{�O��l����ʙ��M��	
�`#U�X�R��/b[��p��lc��Qۉ��˛����mc����4!D��9.�����)�Un���Y�Ϟ.(��0�F
�
�e�����S�����`}��H��%:�pU����3*��)5�%���'w���{����.���ndG�����r�0��\A4���Ǆ
$�~�����t̧�Z=拫�ׄ�H�����Eԡ��WX*�=~]�_2'I�'SS6���J��KC��6�ђ���
Ϝ����uF���k-`��D�l�- ���m�#U��M1.��YkLx�rT,�a:��hA�Úڝ$�|II�R�`��}�2L�����N���/\K�s��h�/�4�b��8;�:O�F�á�i�(�wO�,�W�X�\m�X��@�p��;����UR��!$��1�V*k�ap��
�R�b�1��I?*���Z�M�r>8H1e����l�˓�䔀�O��Il-2��c�)B��A��
/� f9�b����W����_��}���A�u�����FQ�N<���D�1�~󡽣���?����:�����?t��/J�~k�4wj+:2�ܴ�Kn��q�x�&�C��җ��_���^O����g���e:���������	P�yQ�aƾ!c�7���X���'ۆ�7\�[Y�61�Dׂ3����e�8È>�V󔋞�f8h�>��M����R���O7.�1}��.�Q%%�� ����H�ֲml����'"Z#(��Ս���i/'�a&t�	���N+��\�9��f�\G��͂9�r~���;u�*<5��ů('��f�Z�������%?�6��"�ÏkhL�<�UP7��"[����:�i�i<����xZ�}����g_�݌����6�^�Nk#����J�M����/�C��
]���T� ��Hզ�'�㈻͏�2�g-�����݉S�c4�?�l�Ur��Kt���r�>A�Ve��:�O[�K��D`��-䉐h�c�Xs"�H�х���awC9�c!��v@�oB��$�>Ȅe�Y�qb,���k�}֍��ϒ�ސ";x���Y������b���ZB>qo3ṁJ�4��!7��S�C�t�6��l������s�Le�喰�(g�3���u?:��Ƒg(����$`���C_��LԪ�@��u�>
��K$���tm��������/�%��9�i�=����嫷8^� ��N�Z
1k���|{0w��eB�m\�����&3���-�"���a㭥��u���lXF�o���u)�=��o����?�Wq u��ѹ�l~%`P��N鸡�}����	�w�
��y�H1,
X K��yR"o}���C1�p9=�yuz^d�z�O@����O1�ˬ���4���V@$���2���� G�z�\�ae��/h�=�#�_���̺��<�;M;^��C	N"�R!�ɹ��մL���6��^���ȰL��;��2]��zH��h��nڲՀ�U�W��g��F�J�������%l�m`�/�[W�d��9-�s�j�����\�����U\'���h�UVT����x��5��r��Bq�>8W�"�Jz|��pN):n'�6k��;��t<��+71\�ڏ�H%�[(nڢɴ:��Xm>3���pW�־��"�N�Y�(�9Yq��\��'�J�_�˜��K0p{������^k�+f�ֿN#���wǂw^��|8Ā$s&�G�M��xZGp��#��S$����Xta��Z�P4�;|��p�Kn���'U�X�#�C��h�o���x����bQ2�v�|8�c��g��f��_U��)��3qU/� 8M�\mL/q
�U�T�|)K�m��M�,��C��o#O,�#�<؟�6(|琳l�0��)��ض��O��q���֮mv��5�O�x�@޳:�%*H�m�*j��2��Ȟ�C�G%��c�(�)�F��O��p��&yU^l��Spk~���ޏ'��7�}y�����Maw<��O�cVPT�x[�Z��A7��p�,c]p7�۲�0����%�Ud
[�m:��3����#>��n�p��m
	&��j-�$f���1����Ҙ�+���@8�T�*[�Y���!,�"	<�����C�z��T4Hc-���a�"@à�Ԓv�1HS̽q��#:�1�X|IOT]�\F�I���Zf^f?�+=��؁�r78��?�3q�P����@**d�� Ý��1;�%]$甂cv���[��n�{��V��H[C@'������P�q�h���P?L`��cR0�AW����g8�����TFW��F7.��p�����=f�eKs]*�4>GJT�
H�V���R�Ѷd�&���4��ep�7l��*k����CN~^	�
��M�+p�0.��O�L]��%%�?X�g�-Ll�BKDz���/F��ڷ�`C*�ya4�8��U���&�ж�-d#��8�7A�S==x��:�S��>���x����C�
+'���"Ҁ%
K�hX����h��&a�ǫX@����x���V��$�,��v �U+�=���R'��
�U���\K/�����#� X4��k\���8��_~[Fb,!
��������6o�<u_�,{W�W� �,��Z��8�\&7���^�K�왜�L�� �6 :vDw;�t��c���ұ��{�V����m��߃z�Q�pvO�5d��NO��m^5u�b��tp�iԲ��W��b�L�E'���:^��f
��)�-�:l��]~���n�Κ����'���S����xl�j�[6{Yth5�k��2*�#����p�j��꫋��!�*.rF�R�tw��t
�v؜w�O~6ӕ"QX
	�]��5�Bfv �<	�U��r(\_?7��z���9*_�����5΅s;��_�\_t��̵�^l"��n�^�����Zퟴ�>��ߢwsd���ޖ��=�Ɂu_! (��s��p�:մ�n���0�5^ez1[E��z�G�gf�7�ݚ�^�re�N�!�!e�>�x��hfW����$�tq�)�ّ}E�xO�!�}ӄ����p�ۅ�(�C�{���5��rgC�uc/�p��]*bW=�5/Mx�p$O��o^N���U��8+G�������>�X��I������~JqטYU��P��,;9��jf�?�c��K���Ь� ���@(�E�jwZX�y��o ̋���sM�u&�G6��ۏ�����e����Q����F�N<�c�vA��l]n���=�����"�"�%�m�@g�+H�� =�!�><'��V��M>I=����Rݔ47a�4�4��P�2������I�d=/H�>,�Ewʆ�4۵^�z�o�U'��o���18�9v�b/	�������,� ��2��cs�����:�>�O%�������e�ڏ�� H�9�u�i�o�]_�?�������ah*��aT�>o�6�Y�B%��+�l4���]��ֈ�{��c��},Ɠ'��MA�4aLV���*��R&;�K?�:ӌޙ<@�W�ѣ�`ܧ�ˆ,qo���K�h�Y�ܠ�#���|L?;��0�/�.�I��w+5F���,�.'[��;H��Db�W˔8l�zm�?�aO�����R����~�U
ؑ�F���8K{XC�PЦ�s�I���˅Ҏ�)Bi���j�~&�2Ġ��
b��t�t@����WE5q��Mȗ�k?�����=7����u��OV0P�D�ER!���|�+���/e(��3�U\<�ŭL����?�`B�dP�$�H?�8XX���sT�Ŝ�uA�ra&�*�NbX�JF�GhU��#}Qd����m؊'�ky�Ё�=z�x�CIrp�LA��/�{�T6S�v�L3"֋Tz:�&��H�^����kd�s�8my��/�9a��d���|�o�U�;I�ረ�W�Em���,��R4�N�>�U��pn\	hr�$�Y��@���@�A�O��q��5��0�?�T�?3�Y�p���f!Wڬ�gn[����<K՘�
�R#��:�*�D:=�'Adg�"�A?�<��I��b#�;a}g4�>?�	y�zh�C|��K��2�<4�f�/D���uG&��q��H�Ί����J�o��S�'SBt�J����ᜥ��E�s5^rC+���P�,�?����$A�X^J%��|�.�P��fI�]�k\xl��3xz	XQ4��M�밭X�K����K��ll�4���EQ���!��H^��:@�2��l_)W��;|{��Z_����\���N��)����"$�_�U�
1O��{�'��-�[1���pU��aT,NG���fPdri���l��O�i��ܳb�Q�3�=/E�F�'nv��UA������N�1���݀=�Kć���O�#�j���"5�͞�ڄ��R�P�	bX	���9�#��a�,9�G�4���ͽ���l�E�ބ�/a�e��5g� c��m�h���*�ҷ��ᬻ��h��L\�G�8t?����M���:�"P����x1�nv��q۸��R|ם�����H0�B4:t@[A�!�^�|2z!i��)T�.��6}���Umn����\S��~N�.I��䁤�S���2�z*l��DIM���H_�qA������ݶ�Ǚ�I{`m>� �� ����prI�KiZ)r�)�.O��,�a+�ϫg�(���g��[���t��K�n�05��:e�1��ʾ��D������/x]	��MC7�1h��v��$M�&dgI��!���̟����S�_��=.U:[_7�7�S�KV[pm��P�{���p�sG���n����!�^���ȁ`�:@�&2*٧>QpKpD�\,�V�Q
v��iZ4t�\��o~mF⾂��u�(jZ�vu�|`bG�vA����f�������XZ��?�D;!ӧe����W�;o�S�|,�y�`�]b��~� ϥ��d��[��c�!cy��5&�7�,B�T֔��}���A���>V�@6v9�}a�(\n��ȳ	=g�dp���~���訣��g�'�Y�G~#����m��K[��*�1d��ﺢ��lf��%�ya�X]��=��FtP�C���bw�$Д�Ŕh����D��e����c�J�6	�v�R�������6\܊��LܷKg�P:V2�+�>&�0�y�@�^s�0 ��2#�yb���&b:�o�&L�J��>oLi̹
n��+U����贺��P��z��'�ܹf��6Q�*Vr�o�i�	@T!�쪠g���%�8���)��@-���o��T��2�>u<�,v�O bZ����1T}���,��'�-�f:
��k�<���$)K��%�� ����G�ޱ���4�{Ƞ����h��ي�U��I�/Y�e3�k_��	�T��D%-�cߋD0�Mh��"���r���svI��a����l���H�� �Arאt�2��Du[1}{xTS�����vƒm����DN;�
B��)��� d�G�,�� �Ҵ�����⮐�"O��u��6B'dv_�S��"=(��y�&��R�܎Bm%\v���6L��j9��"�	���� �n�[nmw2٧�t��^%��-`k��%]������a�� ��&_OK�wd�4H�:�h����#��vL,��		ô	�W�D����0	2��$7�']�2<�Rp2|�	�H�Ij(1�GwG3�B)�8�D;�N����t5���i�S�
�Bs�g�޺�!�Bv�n������>=��m��<X��ܱ�L:\ӗ�?�r}H�?u.�xk*U6�6�@����t��g�k�M�n,�`~��k�(�"�iV�)��V�9�����Ľh��qY�~��$M¡g|i��l��#�$_�T7|z��M��|4�
��j�1��Pci"�}�� 5M|\`9��pU��*��?+==���4�	.c�����ĝ� i��Q�*Hj�#���]��\Ȋ���<�����9��k��/%��=υ_Œ��Z4�3�"eҮ��r�5��E���7G)cQ�l�6�~)�G���L�52�����j��3U��2:Y��Za�.��v��t^Sj�C��z�Ĕ׮�x=n�5W!1 �%\R;S��5�I��'�lA�|��ב0f����*�U��U�aJ��)j?x
���\M�֑;EVƧ0�������)�iu뗥o�Ҳ!��9�!}����Ɔ��qX�Ec?��v�jc�����,�/_�P�l[\4k0 ���a�\Q���ok�R	÷��v��9 ���C˭fҋ}/�مm�I-���=h��h��r�x}D&��I�m=�\��@h����OV��,�����dC�!sJ.�(,�A1�3�{�n��efW%WC3GH���� �^����[=~ �����sqƮ��SA�Bݏ0ג�	y}����c��@x�+�֚�cj�!K���G �(
%w���-���T�����4�3�;�.g4�aOs�x��m�ǐ5��?���C��dS��Ua�nP9��˰����Y��]q�<"-��*�����gH%��*GZ�}[���Z39+���+�it1����Ր����%��lo���H@M$��Q�#�0�����W�<��ů9/WZ,Ur�� �a�ߣ#n�{����r�X��oy[�e���h��{��A����d'&3���:�Oߐ��"����?�4��϶�Z�M�/0��Oh�u��G����
F�K��o�7�Q��l��*�B�Lw=΅q5�g����5\�A��Z�>v�$����5�{����	46�wp�#n�F�0S*�_���>^�%�Y8�M9�i KG=��i9�1�D��Tڲ� �⨖|�/�k|3�Ε<J�+Oh.�v�"k������|��R�P��0�Ut>籠]?��8~ت�?3�EkM䪚��cP�P�o,��I��EH�̴�,�.�n{�-��C�e	<h��d�&�A���^T�On_�?�R{�Gϯ�����Y%j>�������d��F�$���Ncg!x�A%U�Ý�߻Tj���˹CIڱHz��XK�+�$OAsZ��J��H�T�m�1�1����*U�ȴ��w�~���f!nT���r����'�il�F���<�B�P�Q�����I��oFz���b�脿��@wtԑ���\��Î��)��^ڴ�^���0�j�������J	�3�`�'�R�B�ju�~�:	��؇��a��ݘ�o�k� b*��]^hp��G!�t��f\��yG��AO5�Q ���W������K��|?0�p��&jɆ �#��A���x��s!�Z�U��T$а�Qd�F�	�s' ���1��f��ݬ�Nm����߸�lg����2'�،��g%U�bQé�G���7��Y�ƚ����(���+S ���W(*��_���D�w.©R�v����د��S�SR-:���-DA��o��tU1�ݔ5ClRR}p֥ �k��̋�}1�N��&��u���;�V���)w����	E����ݒKJy�2�pJ{�A[�Yn%D]�1\Eɞ��q������_��yKS�V�����ոX�%�vo����.�����q�*�;]�3ë+E�PG)3���zc ���"��ƈ�:p���Ҷ23>n��	H	P�q-u�a��}N�҂)N7���@m�$�	Kk��wɱ�%}ꔦ����L&B�v{b��+��%��(����%�o`h��u9����?������m��DA�4s�m�Ǭ�>��Pͯ����F���x>l���f�f�~�w���㳲dEH�����N�G�b�Nc���[pI>���o�"���h@�^�b��3�+������Io>p{U��$�Þ�z|��Y�o���W��U�lx>K��H��u��<�N�?H�~644Y~�� �X������������%��N�W��ʳa��#��1\����[�o��L����i�p�K��M��qA��+|@a������3��k�>v������� ���_1
3��7���Y�G����őLǽ�3eje1;��/:���a0x��U�%o:�r�f\4N� }.i.q��"�3-arU/��������5[tY��r�>����<
�H����q'�[W���cwy��-����2�����M�)���xQ_�OH-0�,�&� ����9=/J@�t=T��{�u�D[o�z*�N�:�L(NC���4�4[z�M��6$��8��[��6
��%ݚj�Q>��.�����_ܹ�Dy?��x����I^Tۣ�k�Ⴢ�em"X7�7��4�K����~��~�Y"��큋Ŭ�uI�E�������t<�\]ar��V�1�� ��0�㲹���)�`���MZB�j)�н5<�D�|M�����gbR����O�iv�A�.���_)�����jԸ�r�t�����nϵu���+Rz=-)i�;�B��^5��?�h}�^��3�LL�~S������6D4k�)W��"��	�ߧE"������tc����������R��|2��Pr@��ɯ�����~����_�Rw�y���2��1�ҹ=Y;O����d@��]��AQ>�f@*G|?��rP<ȰJ�|�:�dv�n*�3N�]�U^���!6���d�K"�S�9�'>�̚�l�w�%��F[z�椈�(ʊU�D����H�?�y:-�?{$4��"d�Ҝ�Wm�W��F�L̓�p�3��*z�B;�����ڄ�FJ�V�Ȍ7E�j�`Y\%�g������r���7�������0s���+����w���Xl��=S<�U`O=P �Ѭ(-�,�d�f���
������j�;R)���2P���:V��,��8�I;DtQp)���ȲQ�QK\�����iL:^F�5��3K������}J��5���s��g��*7�����V��H���4p������(M�K׏�� ���c?�/-�c���N'Ц"��V��J�ԁ��I�N�/JA2��E
��'���Tu�v�7V��U��E0�p����^o����@�n^̽&fGw<�I�%Nq���2��ʠ��:�_�y�A�����1B7���刅0�P}�@�.�~r�1�q0�4N��H�R1�V��ņ��>��7�U�}�O��<�ɪ��s�]�9NMQ�x���y��S�X����i� t��O}xW���G�+{��_��PY���xة�:�6m8U��ѝ�ڠqka��$;��GBe�_㾢�T�/�/�8~od�!z��o	����a�Ɣ'����X�i�T��rP�9�C��oY<�D%�J�ڵm���r��R��0<���oӵ�Aq��q��crz}��!����zf�Y�Z���k�%���K��$�T�V�A�_>��yY����`,�G�rt�7{�k{��-�%匤.�
�P2�嚃C?�u�R�D"�.l��=��7v�Huw���%��vU��u1(ku=k�_g�nIR�]�������r��t��fb�7�*Ҿ�(�yv[�_�ʾ���N��u��K>}��s�b�z}"�T
����p^G|��Ԩ���5�m�|���;^X|�l�����}vܤR�Í�t?b=O!� S��?�����,bt��ڿF���@�6>]�:���/6~��Sl��p��gs�:������2���n(��yj�x�I~TyF�m�e-��AK�#�#ق�i�Ζ�R� ��e�I�A[	(�b8Ǟ-�/�)N�B���,��aUľ�-���e�*顉!�o�~� <�ܜ�ִ�w�H�� jJ�V����W"7[�$�+&5)Q%����[�P�e(�HU����$4�6�j&lz*��S��1~��S���z#�uF��K�'_Wo"1��pz8�������^ۻ��O�����z�0I�c���R���m��5w��L!%�xD��Bb�۽��1��Ə<�H4U�3��VP���?=��G�,\�0��a&����@���8�EH���|-N�ŏUmK7}�X�3|��z0�!1?��8m^�i����zJ�H�n4�z��I �f�(�D{;��ơ�ڋq��V�{�MD�\���݈G�<Z�c��JҬczU�*��'��U}�1Ҥ��
���,�W$��>8'���U�UG~�gD�p�k�c�v���+5��хN����uQNp���&�7����y��a�!�ĩ��,��v �0�y"~Gn"��҄d��k>É1\���!c���U
�k���gw-6��ŝ��g��+�a��$m�W?��1J�*����pvB�����1�FJ:e
E��j����-�ӹ|Q���پ���X����cKՑ ��ΚH�M!�]�)��c/���<�8G��|,	s���	9�s��&(}��g�Eؚ-�#�e�i,��K��j���\�*縰?����Xzk.��r���t��� �n�����Ȭ�(�(K��� �2��^$F���H�Tf��gS�3#6�]��(����k��gn򻹶�ƍ�M#O�2-l�enw�o���jS�;�I��DIP!�e���q�ܱ�gw�g��\B<~��X�HX��d �)@8��5�����a�]�� �ց������aǵ���*�f~��Cya�<{�N=q�j|��]�vB@<�K���ɺ��Y�L����?D{J�o쭲�9��0�6�O��n!�2=U#�E�u�DN�)��/&�z��,@l�ćVB���U%�8m4�Xt&)��.�}@�	�Q�����gk��[B���Ƶ,�ّ��	6w/�Q���R_ޡ}���_רAT�T����M4ztw!�4C�:�.b��!q���S���R@�虐#Ԋ��R��O/�w�����9����`���n�콡j��+E��l�	�4$ r��W���Sx>�P��w�.t���{��z��u*��v)�*�xO='^�98
<��{:σ4�)|n��>��5��WLp�_�ܗ�8e��AT��I[�6}P������� ��`+ ���&�h�hy����|l�T۔}2(e�he�a�=$jn�4���'�6�N��,����r��������y2�]�D6Q�g&	Y#��S�&QA�����9X�-Mn?���`}��A�C�'��5("7l�%��Ʀn��˳C�F��љy��˟�~}�ɐ57)��@�^xK]�x�6�UH�a��U�s��)����7|2�TVi��ݢa�y�j���j���ږ	t�����S�~�ҤQ��@������<���A����_�K=j�b����Bi�l�t�r5~x�y����)a��O�h���+�_ڸ�Eha5�w����<e�A�t&q2�/Q���(�P�ߙ���W��W"������k�a�ވ�NS,0���}0!}0�{��&3�A�
j��Թ�`�@R5*��u�k=*�h7����E�Ӡ��l��ME0��}��
�CT��x19�"��C�TOY��v�9�2		]� $��S��m��=鉔�<�ā����=���������K��d<W[��'����Ӿ�s���V�����8�+��K�+�kk�q�Jlty��3u���`�t����Y��v�MN	�О���a�B��=eЈ�oLo-J����_��j��m)�ݧm�V�=�"���#0B��A~j<�=���Xp~�+*v�[�Ya����G�3y��$�	��5�1G�s�?8t���C��ۙe ��ӏ��-Id|�a��pѓW6�6�t!��e���X�-����eL�;�/ހ�[����z������X�L��^�F�.I�I(��6�+���.�[���Yr��!qύw>���D{-A���| �(�uW�#��ܾ��	a;W�N���Eš4�.����2�ʼ���︭�vNJel�=��{Dtѵ�����D$�b4C�*�{!�Q�Y���eK�j��/���ӡ����i�3^���h�#z�5g`R��4�<�e�k���=��'FFui��ddCM�`�Ջ�)&�s��ga�4T7z��������~�)��|���{n�{dE���RuE�w� ����2����!����xt�(��eb�jo���P&�]��=�����֒&��yAٰ�B���ۗmx��K��<?��Q��0HG�#{
�%t��R��P��昛#�j�h��0蟍[���ջ�?�:N�&���Q4.Y72�5'�J^ʃ�$�j%��B��>��eO��{��@����]N�ze�ߛ��M	�s��Ư�O���z]���)�X����s �����%�DȢKu?$p��}gr�Ӕ���!�R�����H��3�F�<�F��g�.�>���G�ZpƬ��uB1GzC�BV�T����<�����΄d��j�d���HV�D�K}T~�$�S���h�N)��B���e~�:z@�w��oG>�r�$��2���m�b��HCt2�Vx6A��[a���v���<N'���n@mo�c�����Wj��`c�TM*Z ֱ����(�+�y�����Ti����&bXxc�8U�[=���/��w����$��Et��!��w��5p49nӋ�4'2Yq]�)g�ʗ�|�����a��s$_nhj�h���'/�K��CP�[ ��#'�Qw��mP~��trO���4�?�#��3��|��HOq��e3��ڇ��7�c�hh��;��t��BYb�ZL�V�?jXy���9�$R �-��m� ��{�D����?�50{���~��!Y��|@�ra�/��jh*�;!�jڐ�r"��q�����+7d�=
z 8t�G���d#��z5��`�8�K�4�6S�%�I<HB�(W����M3����Up4��ǥ4u���J�Lyw����� �[��}��ʑ��I�����$�]Q٪cu�ǲ��)4���-JS�Q��n ���������e�[�&g�4��ϋ��&�����v��@�r��7���W:�,-���ϗ�j �b%� 6�ƠG�l�j`f�fV�W�[��&+c���J���hU�k"����(�Wu�i:S3�'ib��2���k���Q��M��H:os��lz�l��E�Fa�+/�?��5G�<��~�I���`(̗�e�L��5��,�㉩[�N#�:)�����=V��E��J����>��`��1d�B�Q�Pa��+xǬ�X�S.֜1��9;=��z�$&Vd��%F�<
@"_eX9/�C�:���Z!U��nzG�U݈$�xqbn�l�����!U�+�E�b��f�o�a�P~xD��>��1�Si��D˲��{���"�"^4 [k�&��"��>s��&iހ;��LFte��$�B�4p��8����^��-�j�~��ΦLА�Č?�Z���F� 5^�x֞�C�d��C+��	2��zVޟ4�*b#)`�*���j��F̤�
�hwxz�:{9_��zďF��`�y��z��kJ$eG��Z�^��?O���g�a͔:]����Ե�׊
��!��k��x�G;���@fv���>�wOF�f~�HO�?B6�Z�̗��J|K��e�4O֓�Y5���5bf���n����	��D��J\钙SB�ExG.��y��'�Lbeߦ����:����~櫩��]Y�OtF��?5��_iF��g�'d.��;GV��Tz�؞E�X�~�Z)��j�w���Ug?��ç�6P��H�d=Qyk��73��Ө�5��%��i�B��^Օ�ں�%j0$v|���	�x�}����B�-8�~��9�𷿃�7�`���l��y5l�K�\Oe�"#��i���7�_{D���a,%���iD0I�q���	�XLo��>�H����_M���:�-Y"? ' 0g}p��U6d����j�/��+�MT��}�������$[�[M.�i��m�b�/͞�ԅ�
ʕ)k�o�F����5Г��RU��L�B��uS�8��bE7��JA!��'�!s}O�a��I\O�����+�Ӛ`b���������M�"P=�P#�x�Q(s�궢n=�Ǧ��w��z
#=h����G�<t�x��ɉ��8NS����1PZ�%���?��?�Py5��,�|9���o�(��\��=�-�\Y���8�� �<��S�7�����=�@\�R�\Y�Gh��/��u� �.��w��-Z)�
�ҫfC]��MR	� I�5|h,�B�A��׷#��%�Q�B���k:e��eg�ݦ�\B��;��*�	�T�u�zL��Z�$�xc���'{ku�4����(�E_�l�<Ī�������\�o�g�E]|�Fv�00�f%OPg������V�%����W��:���k�QH���|�����������#'t�@���r�ޣ��9n�bf$�?/2b�Q�(ugGS]E�VJ�dݗ���IY6b��#�=w�g��6���wu�{q�"��lo8S��+NE\�&��u���~TS-��մ T=����i��9�=�0�N�(!0��(������ e�mPUʏ5@Q|SBR'A"d@��k"6�rW�vv�+'QA��K�_G|����b��6�?T�qm?)p��#�ABI���78���� P�#}�[�k��x�q���@�wI����lf�	R/h����>
�<D���Fg�h{�u�,}�}�|_��t|~��1D$��}�R��!�kx�h�G� ����Ŗ��scs�E��ֳ����s��N�\0�q:6N-<��.a����4o|*��x>J�w�z��$d9�e�L��A\0�"�%D��~h���fhT�c������!J�'X��G�P�d�\g���]�pNN��I�S̞c srGQ���Y��;�!��Mq%������f�'NYI�sߤx�~��.��+�Q��^�s���ne~A7�s��`% �o�Mj��X%|�EQ[�7 ��)W@�X�}�e�����vq��IQ{A��nȰj)�v�Dr&y~p"h}T�H]eO/ؐ	6����ݵ� $
�B64g�焋���XR�̋��f���1l�4��2;� t!�w#b�N�͊@=Ӕ��t<���8N��4ѿ���FE��k�4��AQ�!�\ߌ:
��J��3���xCܞ�1�fO��x�֕�˳���4͖k�m��4QW�sn�C�J<���H�ԯ�GH?���,f" ,�}��8�QO�ڽi��W���ܦ%�g,�͡+)�	�Eݑ�D�X��%n��҈���~jQ��s��.�9^�:�b�E�$��\Gqح��˭	/�Qw�+�/���r]�cm�ա8ׂnL�RS��3����X<"���	O�ٺ�\�c�Ɯ��������b]F�\&%ϝ1�8���������q"e�_&��m~���͸pcV��k���+Db~�<��NPd4X�x��΅l\ߨ���f½A�k��D�(6\�ч�~�}F�Eɫ�fwQ��+,vtmVa9a�0���,�σ)���m��ŧl�i�`��r�!�*_���J}���Β�cV8q����csX	�`qK�h<�v���y��m��L�z���J�m�>\��^hz77xAh9(#��f/W�?����؆��f�h#F�m�<k������)�{WK�a��\�(H�Meݾ
��e��T* �E�Mw(�*M#F>�dwr�_ذ���`�Iԩ�=�߫��4�2�;x��t�x�� �?.�mA�Q��)v
�87˻�B`��
s�����c0��.�,8O���I�
�	 ��ÿ�U:/�Yp [�qc���h��y�}o�,����!�%�����j�>����N�X�tꓓ�e��WS��e{GGF���`H^���xp|�x`�nQΩ6�|�)��!���<Q�= �o�4ߒ�����C�b�$�>�S���y �-bf�=��2��;S�n�ƴƑ@� ���܆gdtL"�O_�'A��6���HM�"���K�}�ϋ�eBrӺ�f��_r���Y�IΪ(�.₃"u������)��l�j��Ǖ3�&�-�ǆw��:C�
�������& �r��ʿ�"	�u��9�(�Ӻ��#��C�:���p�{;�h�61)���!~�H�$��~���J���74�n�s�%�o����m�y|��7H����|W����j���˷\��1$�m��
-��\*y�lc�>��aRz�P̩	.�3C,�fX/�3�_ֶM�h/�J�N�ך0�uS������/��������!t����{�����y�� ?7bu ��12Kly�'W.Ĉ��i���q�����$����D;���Y�A�7 $%4
e�s��4"+���J�Kh}@�M�����aH����jX��VM���ԏݒ؋���3��]�|�@	Z��A�j <�aĈ� ~F���X��U	��or� ��_�~��'?Z�7�1PU�ЏZ��^�Աӊ*���	�賫p`1��%��}����Kz���K ��D;g@�W«�frei�"�Dq��;�;�E��B�Mr	���Q��AM	@<r��_��:;�@�Z�8!w��h{ok3,�8�*������SL�&(s���Oh}5�f֖�SS͌�1X�"����΄S�fn̐�j�Y��C��Ɂ�>NA˝���;��c��w�"��Qm�_g���?�ĝk�FK��p�u�.	��q��Fv�6,��!�f��F���A��2䷂��Y	�5�T��t<���d�2l]p�`����D>�L����f�F�1�|8��?��WA��>|�2�_�M,�d�(@��R�D��� G}%�1,�nn',���\	���Dϰ��.�|���c����r��>���1pϴ�;ږ�ĠA-`�X	��E*5���x���u���Ds^'N�!(��i��v��u*؁�{+�ʚ~[��6M2 ��?p&�95ᐆ?���b.Q-�ƨlG����[��l�3���	���g�|�����i���w��\�:�h�xX��_�Gl\��
X��̐�	^�ѷ�ɠ����A��1�/�u�p��-MZ'�	.��|%�G����*�g6�!�kl5W���� �ٜ����ɰ\��'(�[ @ZZ���d���0*���˾^I�7S�
�$l��9v�,��-ד��;lT1��_P�����Oc&�%(t.2s;%{�5'�{�����d�ŅYD��'2��K�Oz��"$Pq�� 
Y��57R-���un}c���lm)����Iq��xۖ�fe��a5HP6��U���-sQN��ۙ���-����JÉ�Ҳ�yK�q�@p��c�{z��$��/�}�ag�����R�QD�}r��IV�
�;$�W��"+��
Bk�U��*©�@��@��GYQ����zoD �Us�@4�4UA�yN������~z�]8=d*"jo�g�q<�*�jЖ2bo��`�cy5Ǉ?\
�$���
��)ѐy#�f��J�&���cNR���f�̓�wH)���؆ӰC�Aq�ӎI�T��q�p�)7L1�!2%k��6Y�Б��6�fgt�(���X^��Ԋ]�≟�[?1� ����l>|hA��q��|$�NpA*��m0v'ŁΖ��br�5īdZ���M�CO�P���fT���{��M6�
$Dh�sR�o�L_<d����R�k�Pr������z�~��������O҄�`C���kJ�/`;�!��{�O^�X���ߋ�貢|���)����y`X���#�z���0��x�� 2����Inz�_���57��L;�ڟ� ����
O0V
�lP�!-��?PT��/��b+�'��ē��x��)|A�U�I��v����g���,Y27��^!��ȍ�<��|b�"g&�,�T �-��E�K1j�04-��@�K����f��R-vd�EyyIF�ѩ*�R��L�>�?눩�k��D��ߍ��,�6z����X�~���D;]\%������%o"��]=��:��s&��_L/��=a1X�Fx��(='�Ż��`��������Kf�3;�Q؃����|�￙|>�O�)J���s3�d5��;p�Jc���5:�`E̼���o�hLSG9�
"�*�B#��C`��J��t*��ӡ!�e�W$�33���~ ~Qz���[?�����3��$�8b���2�Hu6��P?R�W�썛��
�4�%-��z�c��v	�1�Y�iP.Hp�6�x:�R����ݒ�A.B�3XB�{vTc>�ıif�
�
D�1,J��}��-���H� �*�ӟsKʫ P�_��!�W>`!WQ��z5��������H�i�o��ɾ`�-i�>A���WtM�o'C�ۛ�7�E)�r(�.�������͑�!�TAm(��^=bA+B"�j3��iv��mUL+%�4�맺�e�Z�ܰ����F��ˊ���z�c�}tpe=� ?�*��]﫫�۰7�1������Y:�N�?�@�:^B-Q�����+'�9�+��[\��-�2ӝ�m��&w_��D#�H��T��k�P������>���;6r$�r���F�گy"d2��1�ߘ�4�'�Od�3R0	�U�w�&�)�@�j�a^ט�^�e�-���8�����ArɈAb��,��+��ZM��A+pc]^�.YN�߬F���#@MX�	vhl@ Nxvi�����^�(�ih��LT��>��^����п�-�d�@<iT�F	�WЅ<�J�����ك�Qi�ll+>���>7vI�Y��Wۆ9����7���C?p�檨W5GuO��m�6��45�c�`��&�R#��ˑב��닉�U�ȱ-^w;=7ߘv(DLK�\�nkZTg�;/�eo�CƿԄLf܁F�R
�x�W:�*� `)�䇡@ #����?�4����.�dS@8Iز-�� l����j�ʉ�g$<�.h"�����i�l���i��c�ϱeo�F�,�{*[�]�Z:�-��|�9<"��bW�Y���U��R���щi
Ty���Q����yQ���>4��狃�O*t����-,u"��J6�k�*�e3�t����[�-�	��tU���Xt������5�]�N�Y��!Q+��ȱ�������(J.�0�꡷�ХM�RrS�r�I�n�t�q5y�V�c�����2G
�.'�lkϢ|7`�W�C#���b�*Y� Yo+��0z�H.V[�ltI����~$r���ɠ���=1�6��}�����+���߸k����a݌y"� ��RA�K�Q��"XǠ�T\ �@��Bp���{X�e���~H�7��?�ފW}R�z|��?s�!:z�DaE��#��������G\G-
�3�ɲ��y9:���5�I�˙���>LE,t��2��~�6VI�&^F��?��R��
Voq7�I�N�a�Z!M�;b&���̫��<q��pq��ƍEZࢗ�y��4u,�F}�זa/7����o���#z��FS���hW��xٕ#=F�sf�,��+�L"���	T��n����R;��c�����T�}eqg��Q�ѬŞ���Q3��8y7*f6?Šh��&��#Ҿ�cp�C\0���`�
Q��jx���@,���:�ʮ�@l��XFU�[�P�Nu��� �"�A""��	�a���J,�Y�ʁ�ՙ+���a2\��o�v��ws�4n�:�=Z+F �}���`?lUi
�\���ê�Xc����?-R�9���GӔ�-�B�E_��ݿ�>���v�C�/�T�Ǉ_�z��핤V�GeV�q���"(L}��Qs"�����pҭ>_ԏ��RY�[`�>z6�?+{�K-��D]ս[�&^|��ē�n��N�Q���X����.�B��]~ō�Ը�0ǲ�V���l+�r;����� �F!�i����R�6��)�L�����ӂR;dڭ{Ku��	D ���ض؊oj���m��a���&u�Й)g�?��N	���F��a�G/��d:���Wr�0
���2R!�����u��ː�z��B��x�!�j�?#mBp7�ʝ��F���c8�
�0ʦ��	4=e�!IRC�|LQ�/wQ�M(0s�E5@��+�]q�G��d�U���1�����9�LWk<���nwk���3�_��v+L}$:��C�^[��ʷt�B�{2��*���:��p���>�+��J�]V�e��Vn:�qu��cc���S	���9��3�Y|z��]_rV#�ky�%���A�J4�`�������H���[~��jz��^�Y��g��@'��З8K&��Wxvh�:2��	=���	�lr�9'�;�-�3�LNRsJ/5�d���8��t5��h�ÚV0d�e
��<�vf���ES�
ËY��_p�WOM�5���I5N�K�˥�3��Ϝ��We��W+<ѼT�@M�h�R�#0��FB7���L��R8n;��|�Z�F(XD�K����6B.��<��6 �>��!*���@c�V�V��.v�P i��PF{4f���0
1 V4��9 �����c���9���W[���H�VB�?9��7��o��y�Sŧ�*��@�Q`����{���'>��d5�-R<��yK>o�� �k���vЕǡ�f�
kŴ<x0��ޗj�lr/X��2b�5�R*�(��*��k���f�X�fq怢N�<0�ҭ(�Kñ��[*ǝu���H���ΰ�K:H���JMB%[l�S�J��T�`�����u�W	�C�(�TW{�Xd/ҭ�k��^$ߧ���a�1!"�K�<_�B�!f����ܥ����v��
𾝩�k<��lB�Dw�`H�G�P}��>Fs��vz����<����v��K�w8�"�R�PŢ͸�f;fS�}�����|a�ξDe����N��g(f���z�t�l��y�wV�f=ό�:'s	|���	�,I(�%�=�Hy��	�4�/�Ż�Y�l�L�o����H�M�p�`.���O>�sq�XdsԴ]\v�4@Z�	zC�~2Q���4��]:LL���K�hn��[8_����<~�rsIS��jZ%�u�#��)01\mQcOW+I�c�c�A�֪�~X�	7����Hve.���}?H�� �[Eal���8j[�p-��v����ˉQ=h���4X��C"�۟�(��M�ahJ��oi#���)�<�c�?���]�0��D�CFv����Xz������=�+g�ɽ������v�^���}.IK���[�<�<�����d�-,���I���j4����oVzàһem�
���4�5�B�ŷ;c�P���� ��^L��nc�*�$_?�؈�q���LT�v��+3C᧡�<锁eT�O����.���}��	����&�u/��~�������b�����=O�Jn?�R�"�n�<J¥hh�����⊄��6�N��-2�ywx� ��:ȝF,g��>��b��������׸�h�(��,J7��EX�)�7�P��k-Kh�l���֬'�!̨5�!��fC�ػl�o�X�Q��º2�bM^��!!Y�*��0f�yt��v|��QE�|*�5or�4�'�����b�҅�cU��Q<����������0�k59�R1<��Hj��*:hqA�!j �b"��А��+�W&�2�2s���R��j��gFRaJ٣8�d�%��Ύ�bC鐖����="%�����`9� ��z+��fd��d0�9l��Yے)��
��\�� 1k��+�� ,�Y�ߌ g��5Xtɬ��ی�p�!G��!}TsB&ȣ���"iN Z�ek[�&�"u�(Tk�3z7�mgN��o�x�qX񳃆�@�f_�ۨ�e&(uti`s��3�M#{�B����*�p��4�1!�$��XFݸ�R��I�ĵ��g�r����=��#2d��!�k۟e�f]��G���axX��M�=o��o`��o�-R���m,��FHF�ut��rU��:;��l%��*ZΗ=n�9X]�f� H��~�wU�2L�/�� +�O�Ѳ����2����r&�
p��)#�������ñ�ԇ��A�J�X�6�K% �-����R�p��Y�*!C�4��)Y�p-�}�6����r���_���sV-*�7 �Rv�	.[sz�;�|TV�y�)d@�{��~ҔVFG ���U'�0���R֎�jt¢%���R�2�5�s���o�R�{�A���a���v� .�J!�qmWq�Tb��)D��gՅ������9�0�_����*��@�� ���㵖�� m��U�*7�3Y����Q�X�ֆ�|��){֭����M���p� �3��FmN�򞢅(�6ba@s�h'gg������ݾ���4��@�����s�?&˸@�<�ƍi��,E���,0�?#�:Ǌ��#(Vqv�6�@Ӗ���W)�����ShJ ":4�b�"�sO�bm������V��T��/��p���V6Տ���/d��B�Y��S���l����\�کS���%L|�����A�T�zp`����
�4~���1u�A���\r��/0~{��tC[� ODX4��
����X�t�x����V�]������5g;Fh� �.K�}�:f\|�^�FM�(�� �(&��6>��|
��?��aH�M%�q�/#���ODDT�VJ�"yc��DZus=��աȞ`��~�i&v�dV0_N1	�S�@��F�B8D����rO���6�?���HcG��f�h/�&{$�<[�_�SdR9�\�K'h�Κ�Ǖ�H��B �׳�[�G�^t����$H|�������C��
3g�]r�C%3����QXg�G4�Rt�䜃q2*}ǥ���;r5 ^�˖9���N�8�T���3����ܡ��?b�>l9&�xG{��$6:�9�����l��=#���h��!��b\>ڂt�.����4\P�a��9��@�H�N�;��'���
��t������#B�Z3Y�aү�+�[�P��F�9��4���UD9<u]J��E�b����Ƥ�� �������n�d9��3�7��̨�֦����S�+�Ho�Z�ċ�$�C�,���2��4�F3*u.FP'�Z�(Op�h2�b|l����h�ꫴlUCr%�6��D$BT>s��������Ղ�Nі���orb��{�:+�@!Φ =�=T�F�vxJ[����ĀQjFɚ8!��&�c��ƣv^&�|�%����۷�Zo+L����hI�5��<�9	8�_ޑ�! jj�yp��SRV$r���h>#�.�Tv-��Z%����P֝^�����jT�>���2��}�|
VB7��dj����T��ߩ薝G�a����w#�e־#�]څ�}�DE�.��^������Yr=F�T�D0V�?�a���k��J	.Y�IAyt?�*�ײ'�}C�S6�g�IZض��c�fZ��9��4���hP��'���x ��f��n�3��=t��╗�g|�	ֽ��=��T�״K!����s�6�z�c�]�����d8���#S��]�d��
] �=qԭ9�m�Z��k_�ާ
Om(�@>�%{���rwj�tE��[[=�>�6E�d}�}6�fWAr��8'�	����d���9�}*Y)ݰ�W���F��5ێ-����ߺ(���䀒ye�x�#̒�f�V�$~o~��o¬���9�G���O��m?8�g�3��c��I�;g�EI��j�3��zG���ޚ�{�XE�]EEj�LXl0�X}��	��t�{�1�Ǐ��#����K�r��h�%_�Rer"��(��U
!�,����(���ܫ<��S��i2,P��YJ]��׼��,��$��>�۔�t�.{��O[�C�����4Rg�Ǜ/� (aUT� K%�'�M�;������ub�~6�g���_��)�[#jfś`?o6���驙�[���j:d�T�P�j��7:�v[�9C�S��*�u0̖-4D�_B"G�\�W�"�v�=�?$s�����X}0���5Kv	 �$c��
g� �3%@Dg� -U� ��+�Ҝ��^y5�R�>��We��^����+#@i���&4���\$�K-��|Ѭ�V�)�KW��UKP$��y���ۺ��O�5r~S�������'%�X+�4>��\��sZ�m{��U�uQm���J�N �a~�`��&3��6;���}�]��㡊�&z��'a�#3��p��R��I�i&/�o!�YC��#͊�� �[�n�v���[���Ӿ{�7�7-��(��OSP�_��F�0~>����s�����<���V�z��,h��re��Y��ۙ�Z��JlW+Y������l�F����W^��l.��v*T���i�}\���*8#Vcㆊ�<�_��X�b���L"p�Ӥ��XT�D�[ ���9j�JY/C�I�	&��W�u���j�<����:��m�E�a����|),}C/���P��5Ht���]<#wõ�ߤGB�B�l������FYը�ԣ�yY
$��O��:"�o�F�c�9N�F�� ��$�P����l�w�j
�{�������,Wb��B����jq9ꮧm�(���֛�D�x���nd�:OuO�p�
����އY_P��ř�3>��9�SNM�n�f��{fY��$SE����.�u$��oRf��ꨏ��S�o|o~�!��X�G�	,K*�vv�˽�VCA���Y�bz"�n��ڷ�)�d]�HC�JL|롘;�A�7�j��ơ�:�a� �(蒬��I�cp6�1��x��ꄥ��F�G����TP[�qܗ;^[�f_�o���݅Z���6j�IڀL�%���+�~��'�\)�P)��$�UR N�hY��"�V��T
0�e�a�o�%���>�}��h8�ڶ�M+}������k:���385B/�<d�  ^��ScW&8���<y'(	�J���i]�`�fϷGs�Z���Uv���~��u-��UI` �z�!%��+��j1
08<w���ҁ\D�T�`]�?Q
����΃�����;}���v�"�k�_R���R9_Fm䋝���)Lq��|qt�鎊�h� ��B�	x�)��o˹����%0��wK�i�6��K�W���d��v�v(a�BQSBxLE��YeM��Y1���,Z~���Ņ���H��	��F��n��#���*GZ�����x��F��v�<��,{�َ����i�B���~�. n�	)�Bσ���GR����V�=7�<���6��}�d�Xd{��BS����6�I�`��� oL
�ݐ:0JVz)�i�����7"l�E�>��S90��$����:T{2�-���/��':^*v�5���� ��ԿM	e`��Q���P��2@��8,����:(�!J}�)�kS���BPk��0��իw5C���W�؆�t��Y�{������� �9����+����E��a��P8?���@lտ&�K2�H׿�R:v�B��~t��Q�hF&Ѵ�֙Nl+)�`����!0��P�-�) ��N�ue��2L�[�&%�@�V�I����� ���ľ���œv���A��_�	
}S�F�>d��F�)����d�xI4��0T�G���S"0�7�@�X�X�^�/Y��d�J.��N�Ln�߸�FU��>2��j� �+i5�_���	��&���5���&"BA�tlѳ�i(�`��""J^J~�X���Tj/��x�mt2(H�B�	0r�����e�15�L���m�. $������|r������������2�V��HM
�@�y�7�#dBt�~�hǰű>o�gc)�(H�ͼ{ڱ=�Ҭ�Ӱ�A�b���q���Z������C��h��G�%�/p��1֛��,9}�^Җ��$����A?t��p��X_�
�(k�^����`����W�/��aO�ҳ{6F@���jv-��������[̚���2�TY��tNU�;��u���`�9��ʊ�@.{A�Q����i����o��]I�0�������%�!��D�����n�2�F3Ͷ��Z>d�����������?�f�+���ʫ�����H�'��8���5�:Q����o�����i-�|M	����uj��It�"S���W�g��L��}�בG�H��D��Ó:�ī��]�a��R�Ԗ&�-L�h(A[ky�4©����p��Y.�r*�A�76�)��?"5G|:9�4u��.
|��b@���Cn�Ƚ���d�6��@ nfz��,��hs�y:�o��a�R@����|��e�����/$�^w=zU�x����>|%�jh�Y�hte���s-���IB��b�	���	�ď�Y�냒d
R峡���梹�(RU&�\v�%Rz�'���[�$���Q+���=���2��E!�T�(jm�ZO��l�/��͋�:4#s�s7n^A�xLT�L_-%T��3){"%/�]�]�K�ol~A]~���I���<�0���)w�&7V���c������,���]*�/�Ѧ�Ѱ+�ud��
h�ն����t�n*������1�E.�;�ݢB��]-��(Hx_i��tH�������l������Pt���HzmB�J����'�,V�w�OXb���*��m ��H�ɜ���R`�*�]y����CيS���x��#V��Z{���\MO��Y���,�:�/�B��9��4?˧cr�� sV����=��������E�K")�py�N��z����Tb�o��W�B]�g�u9'J�/;���[�34���Q!���T=�hV|�Eٰ;1W����V��J�t�b޺VLb���������1�4L����Zï�l�ѠP�P�}[�lD�h�Y��ƿ���J�U$[W"�{��r�{bKQHH���Fp'�tk���}�W��Bm�|��G\9 _�;���?.2t�_��� ����> �0��[9"B3��
;�T2|�MQeV��Z�ݕh{�W4d�%�Q���~B���Ai�,�������5X:�"��eU����c"a��?p"5*�+�IPbޣ�ѣ���r:���;%²i����$��}v�B��Jk�m��O�t�(n�V�@�e#m�6T�<������kK����88վMb����^�^$�R�<	�ɧx!g��k���.�L�����Vl8�Ν����H�n�� ����3���YE�"��'6�6/��T�瓈�m�~ڸx]Gm#"@����YS����U�E��KA?(V���2�D8���O�R�~5$]R _��0��;\�	<�iTYp9�#�K�����k2�����J�>:V�6�݋M32��\&�vn0H�}ج3f�m�A!�'��Ӑl�g��Sx�K���%�̯������,�%�q�z1�+�#%���.kF��ǽ3�wI%Z!m2-֞�Ͼ��	����z�ǘUt�C��,l�����y'.��q���eM���Rފt	�GU�B�+� �P�*?Qʺdb���\v����܍�w���7�������/@���^&;W~�����z��C�gP�i]�N^Q]z�ܪJF�Qd9|8~��g8�⯕_	,f�TC��y�U��lۺmlI��#�8���e�*�gD��Z���z}_"�Yr�$y�6��8��l���c���`2d~�鱼�}�)�@�L3#�'��6Z���F�\+�	��<�["FΓ�&2$ȣ��Ɣ�*���$#'����(�Q`N��Mɭ�O�iP�L��ӅQ��83)#���ҭ� �z�.b?��s����4SHE�i	�� ��0�t��E~0R��2�5��Vʥ���=�X���JW���v�L�dciC�k�$�C��M}�N4|��� R�]�{�ElP�rdʱ�U�\��+��L��M��G��Yl��
�SĿ?���·"/w����7��g�^.0WgG+5�\C,��bwȽ��p�.C�<R
>K���؜L����qX ��'���aR#���t������C*�1���a��B�ˋ��q��Țg�͞J�`�'h�Q�}���$Κ�zB�O�/U���GYm��|��^(��L�����f�e��4����5?�"Qa�	/������K�{���8hz�V���-�h�H���Mt�����
�uc�����R*���Ҟ�vŗ����'Mt@1�\@�?����Go�JWq�l�:�}�Uv�*m��RU6����g���b3�eOݪz�:��(���^�({�Lp3�4����ݬ�Wj��n0��U���$1><ю(�d�6��:�+M����/d�ca?����̷%�<l�D(�!@��+���ur"j��:}��P<���O�=I��X4��Ҍn?�A�e���ct{"���yܱ���s�Ihoy>����@��¦�ϵxs���֜��Ӝ��[O/�J���1��P� �7�%�z`��fRIʵ=u��M)��&��_]�1�j� ���XK�	˪+�h'=�a�1/��{�z{��ȹS�Gj�"�!ٱDy\|n~�<�83����"f�]Q�?���A�#ؤ�[V��� "	C�G�0L�!��mj����K�-j0����j����@$�S�����F�YˊQ�)��X�[�Ȁ
ZL|�!ZP[�b�����.�֕�Lu;���jN�PP�%�}�	y�e���tmUZ�<�J�Ӑ��ޒY;��>ju>�}��z���v�<�I�I+s�$�u
��Vm{�hxk�0��I�!�v^I�'���1�X8������s��Isk���x�|�|���9M4s������W�&Tj�:���k�sz�w��zwYT����du7�ҝش|��n/#�5��?*"�`����*�_e�;�q�S�N��0�?��M��|*�� �~�0���<�isp]_f-n2�
S�g2�S� ��l�=cFyS�]���^EZ^Z��jd�Uh�)E�����}FR\�l�<���hi��R~��*,\f��,�dD�e���e��=��n�������KHT��ԙQ�� ��_5�L�'Ԝ��GؗJ�6Hx�5���$��>�9��g��`����K &7Ԡ�Tz���]3�~,��cs�z���V��Gz@ �V��?�����z(#`Hw���D!�P����+Z���E��HO���u�����""��*Tɶ_��%��<���(N�Uw�Ņ
Qi�v��X�п��0ݧ�ukv�]��<�*c���>�K�|y#m�&x���d�+"�f�{��)��[U��zs��o��]ִ!����M�Ջܗ�v��Gז1`e4��2���lZ�W3�l��7�ܵk��&k0�C�W"#x͢�aJ��`���8muo����D�b!䅒��>�0���`�*�vQ���H}�����?Q؆�*���f� g�?Y��K3뷭�!����%�M�ǽD�FۯY��(e�E�`���8�������o(��mw��ra8� .�\.q�LB˖/.�����n�f&_�O�Qkz����d�/l�zA^�5�T@��`ܦ����v- ��=@�pr[̭��@�� (���Y"���	�16>%;6��_����̍�N!a=�?EK���Bu�v�Pzzݷ�Wk�GV�sXs��!��G�j��B��^��UaZ�)`���g���Ƚ���c�̲��r�G"��fKS�����OH�n�c����[��He�����������y�9�`sN0�7Q�4���7�St�'lw+�DÑ����^��/"%��-*���O���6D�`<��31]��)�Iuc|[��)H�K����!�վ�Qμ�M�槖��S`�M�S�.~�H��PHIȃ��f�7:���t$ �q�s�*�d�o-���8?�Y2ꦕ�p�������4������L޼ń��h�Ko���NL���r#�'� �8x��Y=l����B9_��,^��A��Ɓ5XU����z�MP\@��H�^�\��f��ߪF����Y1�)p*�_��@��|ձ @�;������w����"b��Zf��艳`�sA5��ᷘ����C�L�9�h��N�6->�;�	C�Y�k��W��[����(��S�V�^Fɱ�^@�""u�H�x��'����P�n�S�).Ǡ�g;��Фk7�p�@�]ԫ��],��t�\U��?'1#�������z���i���[�l��Cr��T�Ak�l4�|"�+U�D����n/�r�dHx(j_�4��E��L̝a�%<w�[���#ޘI%��L.�?�Z�Jg�x�\�B�f۫��k�,M�( Bi�����@��Ÿk}��Emܩ�6���d%�{Ю'o��?: ꑫ~"�Ēe
���{�'��#4B_����R��r��9�|��6�o)��J�ww!E�>.�d�gx�?�>;�x�nl���02�9g���Fw�8��*��x�7�}�o�S�� �OܓZ�B-+G����c�z���L#-���`
]-�{`$ZEi�N���^y(�h���)��5Ɵ`���2��ة���ޢQ,ZV��T��β$|�����O��`E���Ϝ~X��Y0iN�������R$V��t=��#�3��*��7����4((�� ��ǧbz?:��	"v�q5db�����ȴ�9�^��6Ծ�{;�(�\�+�,e��122���
S�d�L^v�trn|���9 �
��C3m�/,������D�+�+�������B���Ue��`q/�E���qW&c��B,��̏X��b��%�b=�*5zr��|����	�F��n~T4�޷�9�E�G@^O���~�'���`~�4V�C ����?xC���qŋ�n��eC���2`򬧣���������`��Z�G��SqFm�8-��"�p�u�u!4���)JO�\b��6Ȳ�\��A��Y�拓^���P;��g�8i�x�%
���j(A�ێ<��]�n��_���D�vt��IX����#9�5�|�(����/'�~.����O��A���_��W�e!t�\w�|�� B�,�����tn
i��nk�E�hI�
�䉂�v���j@�Ԝ�^�)��F��I!~}��Ã��K�q���~� X8����f��lR��;�����V��&�Tt����^~RWۋZ����%�=��8�2����3��+e޻�3�8��h���F��#�b��Dy�9����V���!��9���pI�h~������t�K}K�y���O���/yEQ�	B+������n�ʶQSU� ����p�d����W��Rr�G�	��J�#�x�Y'=0�&gQ��n�;�M+6���� 9W�̌l�H����I��6Z]���p^UO���-]�/U d#R=F�ԇ��2��XРJ�W�aswy�F�G�5H���Ze\��HD�pق�md�á��D��ºJ~
��&�.[����h���h��CD���v9M��n��h��9˔Q�h}��r�E�j'�G�$�N�d��|����#m1y�7�F���	Z>��*��{8��%���
o)n��=�~x��Ůެ9���lw8�%�׼�5��=���Km �f��i4�3�T*�KIe(f�-���6I���<{�lJ���iS���K�GͿo��6_��,0��������1l2g>�3+ǵӀ��Uo�_��Y�ъ���k�ݔ�prIzn�`�@�:�:�	q���v�@��q�#��F���/\��1-b�"��ö�e��Wj�M<�|�qf���@��q��8���O�1�虶�WqF|l��El$v���;q0$�voI�=0��L$�Lv��H1�m���]Ͱ��isW�>A
�;��{�n��F&�k�-L9p�'=^�#�&*	���eu	�����f�=�d�5? ^�`d�=Π�>�_���ࢳ����t9~��|�$��;9WW��'���g�\9,u+�/:y��.�8�)����;�|�:.r�kgY�`�Du������<����� p<��5�k�s�~�*6E�1��4NR���}�cAX��g�Hə���+�7.Xd�k���M�=�dK�%�]*��D���3R����C�軈�>�\TS�j��ԟ��S����3�B�y��og�g��s����0�f��ة)�I�����+q(X9nb+c��k���PՂ�9�˿��������A̸�غ����_����q�U��a�[�Pr��=�Ө�fq���:F��|.<����.��� �\�����s6�Q*���d;Z�Y�I3����IP2&R�%��}b�8(���?w���+�����3ߤ�Xl��	>(#B���/�?Ԯƾ�L��z�4��]8s:P��|4�f��BdXP #�7��*ܴ��ǧO�*�G'�S6L��Z���G"q��̉'6=�E� ����L\��b;*s�҇���`s|�Qn�T�O{e-lEL�f���AW(8\z�6�a_3�_���[\xzTn�ڨ�!�cJ��(�R�5N'�t��c�(f�6>p:]w�Iz6~h|�tR\2/�#0�hD#����vL�uE�BL<��g����o����,4k�Џ��,�é_-��ͼ�Ą������U������h���:.�;]ogv@x���xl�2 E�$5��K+2X�G+`k:��E��	��K��T5�i�'�#%0?��χ�G�vԶF�f�iU���E��XzA�d}����42����֪辎B��C}��d�
�Z�5�zYn�}D��k�ܒ�"����CP�]pLؗL99n(Ɯ�Tk*���%̄f>e�29 J7	�LST�zcp���\�j�VǷd�:e�Oi�>��56>=s{27gП4�c}eg;��}CEi[}E�e�)oӃ���8����Oq�X��@�y�����[��� Nhnx��ol�Ϭ��qk� ��R�#P��Z���U⓼#/��'�S���P����a��́pԌva���3��ZU9���*����>~��`{K_�&�zA"�ЏɁ��s�NO�\�7�'ꀸqj�z�O�Η���H�Ј�Aݚ���{	1��x^�V���v�@Z��:���*E���>���K���r�_�qH��"EE1թȕpc��>��D����d���`'=��}<��z9�a��a�A݆�O��bq�=���a���Ņ3 ��W���!���<'/hQ�j �ǧ95�e`n^T}U&�0�+��d����m��'��
x U��k�L]��n+�:m'�&JS�Wř�=tD���?�]���d��}�� Rv������/p>�Vzn��a�w������&��`y@l�Y����}	>x��J��� ;�U�X x{�Ra�Q>�QAK�+r������B!D�D�~,�^�i�'�����Fz>ֹGo��\yM%�����4X��Kkz[Qآ �����vUۛZ�8ڷė�Q$���H�@ոQ�G���^Be�LX�����]�'�/��S�����u��d�l;9}��~���K]x�i��Bc쟞ϗ[4='o�Y>0�R�@�3A)���ʤ`Z��V_� �IZ'�1Q��!��8�nwiP��v�p�t�L���r,EQcz������Aeq���P��~�2�(�����C#�~��D�'-� �H�'<U_��Qܨ�9�`�+z�+�����|�����ܽ+�ٛ-�J,��ˢ�'4UA���5��t��\����L}TI�v@wN5����m���,g�[g%}�/]��N*e����V��%T$4Wo/߅��ʽ����H2�v�����II����H�'<Ji�q���f�v�f�>'���L额 �+b}�?K��D�,3v��"��*B�`v�����َ_K��2r�C�j�ΚEo�ai7���]c�t�E�|A��:�Mq�I4Z҆E���1&1�^dȣ"��}�	���=�}}�~곁�<��K����#)�L�Vc�Me��v�R ��o�4r.�U�T|��k���S���ψf��]�I����*5�ƾܥ;d���9s'p�v����!�^���VT1ͣW�Fʠh�f��4�A)��\�d3O�Ս?�8��g���}�9�'R���ID���&��?ܕ�G
�?cIUa\�z>���A�A��l
ꂲ_;�"�b
ZR8<���2�&��K(����ˀ᣹hlhe�� %Ơ���K��6r%,��{����Q�4��f�#�^��Lb���a�����3^	������x[��/��۽��0`[��F��U�v4��
L����f $*u��oT1�e�3���=x�Pޝ�q�aA�����Y�2AY���1d��PiC�ދg�(լ��T�i��ȵ����F�'I��������^+�1O��Z��~Zb�cG�� y��Y^i��6fr�g�<�t���~�Xh�z\ϯۭ��@R)pI��Z^���Wx(�ZI��q��f-u�W�0�%��W���Y�����"��nxS����=k�s�����y�P���	�'O,l�0d+�z�N}��E<N��K�V�z�'?S^��K�����V���x�).vu���O?b�W�����w*M��=�4�]��J1��F��a�G���e�p��n<�*�Am/�n���+Q�+#� �_�y[t��|���.9#�4�u�1s"������̲jߍ��z�6k`<��f�GP~~��E~Ψ#��b�S�����Ӛ�/I����>�]��@DF�Kh���n+���[Kd�w9��=s�M��"� �������o%���x��_�5�ڟ�11>�^�M:���"�.��A¯o��sr�j�k,fǭ�5�x��@Ȼ�
ثxa��;Mi��Uz<Inc#�@�*(bĀE>�&6��Jx�j���:~-(^��U��@g!�� �I�
�ݑ"�kJK�m�TڕN��Xv¾�� 4*����$�؝�9`�g����W��/�۵�%R��w����N;j�o��Aw��ȓ֥9B�ŕ��M�%���8D�nkPK����C+�r����l"tHJ��-F��q��*��(I�c�D��
0��h�!��L�4[���(v���zx��Z~�yV��kV�L� ԥ����88���%85M��ǉ�?J�&�hgG>Xk���w#��:7;��r���W���CC�w��s���ǑJr���^���qC��X���L�o@.�R�F;��5)�E��U���d(t�����`�v&��`d0�k��7�9����M��GHjK$�F���z����H�0oȚڈt��8�8�^	:`4�u6d[-��M��l���{k2,B;[�&����(�=*$��OnZ�Z= ���0�}u���� y�F�V��#���t�6��4w���'(�͚�H%�!��8�rFC`1���e���u��ޞu BTܭ&�E���0��<k{Л>j��y��x�_�C� l>l��ȏ��]�C-�VA}���1L>�C|ÂZ(`72�ct#��:�g0��ח��-����� Z�t4�-z��3y4�R$�7k(�TI�ɷ`yL��� �jK.��C}�	J�?���e�Mb��줚|���~�AP��.E��S�&^��mǉ���Gg��n�nD�ʨ<h[Ap��6>�y���R�;Mf܁��D����#��'�ptye+[Gi�S��}���q���m&ln�Lx ?}�.b<U���y<�(���0��oi���j	��/�ߌE�{�b����~�>8m~������4;@�5f�07�S��&\-'�'��\j�=�l�ʀ�w?Y���ߺ)��o�0�����������B�<�9cF�fpZ�P�prQ.(8�����q�3x\�C��6�������Į c&`��R�=L������'��� �2U	��������~�&9A�ڧds�Ӑ-q>���}x��Z؟��H1�8m���G��@^Ϻ8�+|3���xp%��D��նH\��Fy�\n���p�,��H�è��/��|q��B�9-w�w
���|�|�=k�:9����Uh��]\`|R�o%V�@o��m_����ʩ�]�J�������S��7P^G�LǕ��úꨅ�U�7w�x�/�/&�#~ǭ���]H�K��GQ���H4��k;(&��^ο�i�(ĭ:\������]������~NX�����A ��:B󤱘�c�,�i4��.*�h
L��V�~� ��gG��F���M�A�Z�5�y��k�*K�S�����Q�/���S�Nnc6Η+1y\����k�+�<��J_�s�6�A�?�wm^�g>�q��u�'��qį��_z�b��g��y�Z�'ÖѾ�K�)�ƣ�9/z���n'���_�Ư�h��7���Hk~���,,��=���Ɇ��8bx�r���U����V��%'��s[����ڇ1�c�b|MI�3p�t���\m\h�o��z�l�ZJ�w/����/%R��mm퉶K>�nW�x(�(r�u^=��tV]3��%
q��G:��ǎ����j�[/��ٹ:�0���7�o0�"����W�����54j�����`v@��Ȳ��{���o���@o��Jߧ3{d�+�2�w���}1OE���k���L�8��h=�C�'5R�>���ⓞ-h�聼�e�����,=�ޭ9`�������An����o�&_���x|���E%�v
��X���>h&(G2���}^+Eɸ/�-$�8���6ѻ�MGm�Q��zZ��?)�BBJ�+�Ү�����t �[�EI���cz	��SHR�,���3Ư�L�Gk�L�PR�3$���/ s5��[t�䫔ۚ�������m퇌'@W��9�ҷ�i��8�g�#T44���vg�skVl�̫�z}��X",D�*H:f������c��鸤}����,ݝ�$=	�e�'�F~�H����:|J���i�xN��(&���U��g�h�H�X��↭.�Qa�A�I�ֱ�4H��B��a$�~�E�6��U�e1;pt61a[5�G�J�l��*���,���f��c����F%s,)�m^�m��۠b������t�y��Ѓ�a(q���?�vW�O����H�#>��vɟƗ#,?UR)x	��͟D�E�xx�$�)���BәA}QL��A������0CD�C`O�/e�HGurc?�&��ާf�t?��	d�>M�c�1.,�����:��&�A���S#à$�D��_�J�L����/4������;�h�3��k�F��#V��A�B�L����:�)��a݇`�۷Wq0�ZDM�:��Ѐf�*2�a��9~$�F+l4����#�j��b)zM���i�R��%�`�t�<9m�}{y�U8��{�D��F��� :R �v��#�
�y��1"-���n��,��C��h ����4��THZ�e�@�}��8�/q�8O�e鳱CF�h�P.V����#xu���>�D��Lԣ�J�����$�{����'D ��Z(�$5M'+���.�����KNq
\j<��
�p��3��
+�m0$\?k�I�Z_�H�h�=�< ��L�*}��xaA.�M-�8���`�uX���3֨�Kl5��"	�2�9Gv���D��:���ָ�o��GY�$�W]�ǫԡ.rg�eۧ�kP�\i�1�I����=�<��KR�
��~�RDW��V �r��[	�pV���o�������W++`E��{n_q��m̪2���~6��{/J�|�u ?��t�ѥϯ��X����L0(�3H�1��gB<]j�(�	�<	���U���Ƣ $�s�a|i�.�dK�C5�Ҷ��t�1?�)���&'����op�l=[����QV��y�M���B|(ͷ�fL�I��]�3�j��X��Θ���=U_I	�Y�4$q��d����!^b��tţ:�Z6��ar��; %$�	�.����M�W[
<��c�/!���SUƊ�v���L	B�!Vc�W̍M�1-3����]:L1w^��w���ŕ���-��=��o�o�����n&�*}�(t� �j���km��p��tzj".�M��@�0j�m��I>�LOQkVX��ܶ���+�m{Z2w�yJ��i��Eb���,P�/n��.�s��o��y�9��@�|�`XVS�$�r�b|����$r�<)��܄Y�JYU��=�v����Y�#�eg'c)���-k;W^iRn������SQa�k�-�솦A��{4�5Rhz��0~4d��D ������_���vh�2V@g�PP���i�ȥ�0h?���Nda>��*��@.�.�_ނe�qk���C�B��Z-w~a����n\��iv�s��^So)�k�~�r ��*FR%�	g�Rݍ��]���K���\|�"��V[�Ԡ?$��Ӓ�^�w���Р�[c�L��< �rMxƓ�Ά���p�~T+�%3��� �Ӛ�m�7�2���U�e�!_?>S!
��>��'�4�9���O��39g�+�1U�l� ��d��	x����&:s)&yy�ѷ�z� yn��_�n�B0������t�l=0�oA�� ���,�𓨰z�#��x'�3��г ��s�v"���s��i��,'��y@'zz#s3L����p��g-YN\m���8g��zk]�(�T�'<A�nf�-�>�b�K���>i=�fr�O@W���Cz����.�Yw���x#�Sȩx��8K�dR���v�7z��Pq"���e�ݔ��F/ѬZ����:�;�a�KW��M�-�G���<����P���9Ԇ����$K,�������T����}�ù !<�{��x�w�ϭ�Av5J`�����L��~���=�?K?k�/ѐ�	�kGKJ6����;����=�v�q|�8h3M��:����8���k+��Y6�Tg[����	>�k��!��	�҉�_����pf�{�D�x�(+w����qO�j_��Z7���^��h��9l���o�j����*�i�̇,~�&��EƩ&_�e��y^}�"���oѬ{�~�Ş1!6/n������4�p�9f.Q^�F�	9���X���Mh��9 v��W�\	�ᘫ8��Ǔ�q�b��o�/ɾ��M�l�꒡3e�j,���-7+�u�l�AO�3-�L����*i���Lͱ޲p��LU��T�O�k��8�Wj3�%F���E,>J-��T���~�qO��`$�w�����޸���Y_ލ��$;f�.���&ǻIB �F������@�c
��JR�=G����9���S3Ng""�7�,|�à�ȥH|'$�	�W���k������r�Y�a��^.�%� u	?ECHC�� ȱ�(Y9n�:u\L�'��x���on4�q��}����N~���?é��&�c%yZ����-MJ�֔&%��~O^�]�t;�"�^ ̓Ϯ�A=IW&��F=p��b
���������	��wb�/�K<~_(=�&���~�ij7�P��iGhb����C�^�L���ZL��S��#���UP�&|����c��$ �,Ȣ��&�QWQ����9�>1��ٸ(u�R����aw3j��x!,��{��\�T�@��Fl����.BG��~�(^�Q4�nG.xX7X�:���aۘ���t��|�Ѷ�)C�a�׃�,�o�k��`7$���'uEF0_N_vun����4a9J�n6oG.�e���bB*�X�<ׁZ��Z��./�=�{�.��L�.'��Bd�F��&u�-�P�
�뱉xʋÜj&CN��6��o�� ���\�v�n٭�ֱp��&�!'�G�1�&�r�"��%h�(Ye4�	�L���_��]�x{������5�4ˑ�����������H�$�ĈG�#�/�y����Ī�$�����>.JAŹ�]�D:�]#!��M���!�,|�gU�8����B����U٨��6qA�����o\kO�BEҚ��#�;�o�vb�(cC"6�*��T-gv�dt�7� �mt%{�G��TG��,*%�kM�gqb� i�Ќb��Tm��$Fqb�"67z@lĠnΟ�q"�]TԽE�DIP���
�O��o5��&��o��`��pUMQ�RKP���$,O� Yzv-�5L�<�)�`���/f�0��)�3}�1��2�$�ʎu����]8'���<���C��9���3LZ?�B�h�@��>t��ڤ������1}o ����ǡFa ��I��h�/�M	Wы��a��@��p��)��t?ø��>��<�d��9����%�?���fkZ��ސMZLG�XB9�{'���H��6���"�x=9�n7�<g�^	��b�{��������:�W�·^c��x�0�������w6
{=[c���|xybfO�_�v ���3��MD�-�-|���%�uV�Dg%�iO�N`�2�t�0��*bR�S+ۧ, �SCyD�Br��>��&�Uwc4B��N��j�l�Y���ww�����u��ޣ<׆T�2��K�x�a!EGo�(�N����~)~�N-F�?��b�=z��0����רSF'95�1%�֚�����NΚ.2��]��⒅��>%Z>u���FX���t	*�Ɋaip��l����H��������%.a۪Hi$Rlz�5��~�	�슕
!D$l��Ӈ��r�(�rZ�Jn.r?���^�L�vP�%��^�m>�g�A[ke%�����;v���+����E��&����F�U��ex�o퀿N��f�$�N<2��>i��y�SU��_E��s[/ģļ�D/�E(�)ޞ'�H�� F����ђ@��mK��{���Yw��{�-x5{�����Wk��)gF�:�j�-�-���Gsg�Q���;K":�"i!����|���S/�r�>Cd�C8R;��ح.�4^ ��/KgF���_�j�2������gǋ�-�����S8ZV,K��x�[����S��Z�"]D*��'&��X6Sҹ!biC%�!\�a
�/�uX8��D>�jLI�ۂ��x9����<�Y$�m�X*|>��d�.��7�N����+ޥv�{)
�3A�u"D�KF��V���oI{�+�+Aa3*�y ��p9xJ�������D��x��ޚ\o�v�ۦ�N�ظz�ϒ��4��g"����q�I�A���cx@G��� ����m@pڙ��~�\oi��p��`��[�N��K�&ȢN��?f���y>M�F�5�r���ѫ��3�w<�)�/RN�}�)�v��0R�Z���Xm�;��$֊�G�L��e%.�ݝ!E6Rm�R5�:�ޫ�����
Cɔ$<Lt!AM
�d��V@�5�|��^%�J����5��m�D���wQ
�,D�A���2�<v(��]
v��E
�x`����@�a��4 ܉����C8K�M��<M���.�M;|SG69�]e�׽QƯ�!'�#IIQ�e����������z�h�߯f�h���~}������H�P�°\d�/����4فh+c�0�f��^�C�/���k�P#X��&�OqK �\�p�W�W�^�Y��MKK_�Q�T�ªf��$h��a�}� l�R�	x*Y/��A��� 0�X��&�J}\�U	ΪFt	��Ei5�ܝ��=�,uX
0��o2��ntܰ��Q��E��>>`^�M��-�^k���5}0�R�}=�����"d��3@mU�R�zUs�J�'�1��\���X��`���Ҭ�?=��0� �q�A�{*�
��`�bꉤ,���M�P���-� �m�7�(������y����C�d��k%K���& 0NF�W7L{o�jG�r^݈kޒG��P�\A׎*:S~�-�,b~�`9� 8̂KY�ϼ#f9��bvF�7w��Si�&���r��+���oM��Fq;����v��&�u@�����߮���8����jҊ�V �\W}��e�Tzu=�'ZCS7� Լp)\R�s�a�i��G����gD'�S�״��ّ���CN@�-.r�x�l�-���!ڐ�{"+!]{�
-�N�*؆�����z��=u��-+V�6��߀_+�a5MK?���c��wA�0.(
:��#����x����AaJ�&�[��ùgx�#ve|*�T�9���/��U~{Шv�=��0��L��>��&>���DP���h��
o���-S�����f�T/f�,� ;�G1k>L�1�r��~�YA���2�Q��;?��md���*�u|+�PqK��rG~��7�A�+h,��V7=�LX���r�NO7����� �5���|���������y:�U��Gs)D�i�D�}I��m�樏Euu62���E�����J�,��4y=^���)�q��Q/'��6�����ɫ�h�}�lG�l�9�q}t���Xӊ�q* �9�ݼ;��0t��6��o&I���?�P�3�Xi������W���\sJ\�T)�l�_a���`��K��n��=}D4��l�����W�h�I�u~�}	ճ��J�A���qa�?��&Dj#�`����|G��g(iExp�����Ғ~S.1��?ϗ�v�Nb]�e<
�m�rɀ��C�|)X�Z�e="K��!���oL�q�����R�z�g1Zg�`@����_��h}gA�OE�R�@�w��\Y	5S�pYŠ��_I1Gn��N�9�h���ļ�V��j�{W�.�`N�P�[�������F"�R�;>�eN]�M���2m-�K�D�u�/�g��TҔh����A(5�a��O�|/�'�Z�u�g����5��˫g��Ǭmj�4�sW�Xgd���O&袐p{1���e�])3��x�u��
��#&o�L��q�̇�������7�4��k ��IF���^VO�߯xm�XC�| �m��ɀ���a�T� $�,w��qy�9T!j[ޖb5a����"Mu]�Ӟ,�u�x���@n�T�#���U��ZTh$z_�hM/J�~lɌ"��P��措s��F�,�uL"����V_]~�A�j�@�;���D����c/Ѽ.��D�q
3��F�D�󳾈(���#*lq)b��(�6#�W�����`��}Ţ���Q���KB�o����x����#I|��e�LLTh`��;3�)�TH/���ivG�w�I��صF]��z����4Y�����2!�,v��qoTI�8��$��<}1��@��<yRA��G�8�Ӻ;°hܡ�K��t��I3�QQ󚢷0����i9\�Usc���im|y��RŌ5j��g�X������iX`UL����1k����/ݬ���tT�bJ�-����V��R>�i(�x��K;�7��s��{HmҮ'�#�W��8@�]C�y
��	�4JYm����B�ʳ��d����VC�Ɔ3�l����p<[`m��m#�)���R
��{�B���ּ�Ta5D���W���]_]#�8jM�
�0J���]<OW��H�k^�CSuV*_�dc�)呔�okP=��0`#��uuU+.@�o�%Y�錑�y��!7�����]�xq�Cx+����7��s�zfn�x.#�|�����>^�Rf]�y1/b�Z����ܶ� �M�������>�E�(�i$*���������H���e�KKU��G2��T�}�`x!4�����W�n*ݲKF�Ӊ�!|9<�Ds����a��ԅ��Sc�|bϢ�c���e�?;��PO��M�?�s�]ĺ�Ta��_@>�[Un��5)��RD�t^�'�4W-@E*qF��t��!�K|�ɐ�3�	P�t�����q�?Vu� �Ve�hz�0~w5W����`�jNa�2�=9t�;�4��0��fq�9��a�6'��u��|���B��s��>�Ub�K�/��M����./�+T���l�q5�T�8-�d�j.���YO1�ߘ�h� j��僋ihGS�������!�2;�<v��pE���S�x�ν��'��h�\ >�T=%UX�. ��p��T��Q�ΎZQ���6��z̸on"�����L�����RwjM��=Ԁ�A��V�������^�����͂ #�
�:�H�<|�쑼�&,���.�<��q�Qcr�����g�=�M����<�� f9���͠D�,�UT*��K�pժ"唪�u�#�,����S�{r��OO�2)ݸ$V%����ӎ�7�22���W����^��gZ�KX�e�O�f��'��k9pF}(�>T�
u�둳���c�q��M���@�s=�3��R�K|�Wfa�����Iw�Ã�b�,CK{�1V"����h�Tݷ�
�%b�\�P���U+m��+V�P'��nN��v�{�LF����;|�n��Q΄X�,�pz>H݌�����n�n�ݓ�k�11�qz�Ywk`����a9g�X�H@W��}�eLί	������(De� �{�Ɣm�봲���k��V��jdl�� I����`3�$��|x/��Դ�dÚ����&����H��jz���y��� +�eU��F��x�%�����o�+B���z�%zmo>j�$3�\7�ϒ{U=L�S���Hx����gf+/��M��}���5<y���dA�J�ê�P{t�Hݷ�<�5��J$�E���җ�&F=Iֲ�$R|y���yP�r��眲�u���l�����g?pf�9MCy���-b�7l��/i�_��LdL�.c�D1E���&qݢ�0���>Yg�����>* �U5�\B޹Cbp|��%�ڡ\��&��Ct��/��O�ܣ���_gj��ip`63v
֖J��[֋7c��|Q�a���a샤ڤ����$�׊Q!eZ�q�~��&�T42��nQ�3��ƙ���J�9��ԝ�}4~}� �r�p�0���=�(��;y!f�?Q"Q�+�A�A[�X�is�ƅ�����ѭ��$�M[��y�Z)���C�KëB�H+�FT�'*�R|8W��?p,��oo�c��W�?�G'�?�����B�2ۺ6�:Ma��`�Qw��Ww�J�%�zB�7qݶL�����U�=;�(�Ҋ`2��82����z�,�p�%x�>)�h���1���29��Ob�d�n~/Q-R��@4^F�
�3T�0~��y���j�=^���e�Zf��%ɜ�"<@c�<r�|
I �u��&o�/���1�F�P$��ol��#���Sp���!�!l�h���D�8����Z^"���]�Ӽ2z�uef�%��5���<'mJ��|Yk��?G�U65P��M��s�GW_4�?t���-�C��a�"�aGv�V�ǎ�u�p��2���ȐφT�gZU�ٸف�$�e�/3��5Xwș�>	�R����,�`��<fm��������q�[N$3����%�_d��ֳ`�ÛN ���xr9TO��n�o���L� ��	 ��{(����������r/�Z5q�- �I�����jݾ���@�E��@X�v�[���|P�?1Iǥ)����M�����J��Q�q�z�T���8��ϝy(/�V�q*�.�O �-"��mH�����C@�R\	�-|�>?&��[�A��������RU�*�Vd���ջ�	=X�g-vE��,<��ME�œ��R1�~{�P��+3�,�����e�k���]���#W`f5q��=T�t���8H�X�خ�F1&/+�\X����B�Y���E��^+�!rz�/�����h[6 '�4���ur.�	:���(~s�7i���e�LHo�D���	
�"XH�b����k7��ĂZ��vA�1D1Mq�(QϐP�~_h�
�����h�������z*�`c�Z���Gr�d����Έ��Nt`w!����0���VT�<����ӑ?\�� >�=e���{o����ͱ-TM��P7 �4�O���Z��G|9*��0t^F#�E��,4�(༴.4>�5�5N�ll.�!K���_с�;�\Z�S�v~i�p
pN٣"r,���ü�����8G��{��^�N��&�OF��������p����A�D
S?�w,��h+�;��P%c�S� ��S=b�2��gY?�d�;��N�e�)8�ݟ�������"O��u1 ov��T� ��IW��#�/�\��!�ק�d{3~���$ʞ��mv��d�-�q����r� ���q��̷����_�T{��>��ڼr�نf<UVʆ��|W!bW+ZH��Vܨ�q��lD�4C�_-t�\�ͪQK���2���	V)��`RX��}� ����`�nၽ?Gw0M^D�/d�}b� w���z�^Y���ϭ���R1W���,3�SA��m�ּ�k���
�2�X�*���X�ӱ`�<�8ʜ�j��^۸���b���&jV�%s?��B�������ޘE(�575\i��N��t��A.xk"�)
�ٚ�mZ�y�_Ig#�6��n�9�K�$e���ԥ��n��� XB�u��6��hc���l,ZG>���Q����ع���uDce���B�ݕ�/xG*��ٟX�UP�������&-�-���Aw"����� I1�A�H�C�� Av�o)��������ϛ�����|wn^�PY�}ό1D�76���]�K�Dy�zbb)��:Qv�h1�?�U�vV�6,�z}]<;>q��a�?pƈ��f��Z�~&"iS�x��~c��(�����)�.e&�_
�ir������ ��wj�妎���C�KY&��}��v�Z+���H _Y��Y���1
�XM�Y��"�H��C�JmG�W����9n�+;-�w���nUv����qΥ���Çx#�1R]�Sߨ"��[41��-��ʣc�,;'�)�5?!��_B�@��a�N�U�"�D�����s��\/���Wu�U�$��5����f0,uI��Y���O1�%�!Q~��Z��kN:2-�}w��i` o�Mx�������x��oB^���D�Kꓝu������Q�''��u���w��kΗ$�;?8^6S�B�{���qp���������j$.29DqW��C���h�{�r�4�
<솾�O��n)��}�dG���GOx_W�a��D	^`��hJ�j,�������Yn�Y&L1#�vcG�X���~3���U��M�D�$��*â��_�xk���;Rج�e=�܇m�ڟ��q�}4:��(��'w��z�9J@���E����:Kgo!�t��Q�K@�X/��ŕ���4	�e�:-�54�@��O���Nū�C,�E���G6lje������O�Z37��(�:��m�b7���^��."�	�M%��[dx����!�W���P�i���e�,ف�2,��|Ym�F�P�K�A*~��[Dvċ��2ٵ����0��iҩ�_��䪩+��6��ǧ�˽ϚU����NrJ]�6��6)��z)��l�7�E��포�?� ~��o��92�V��_�_UH��*����P`���&��s���IP�A��n�?�qx>^��i�cJ���!EmgٖՄdI(G޳�C��PG���g��h���{���}E�����cg��� A6ghQ
��m-�Z���Е���
)�[5|HN�15M�T,��t�Y	���2��
b#&��!�u8�|��`�݈W��2��'�M/�=�Ŵ�U"�ȶ`|8�Ԃ��6g{���ef/���&�RwEm��(� y�x��!ޯ 6�ϓP��dj!�=��"�"�f�YC��V5�UH���C��֡���?��}	�|ng˩�]NĜ����T�	۪];~U���>W2D��:�'z�IZd�ʛ�u��z�/��,�X���_��ad�r��ĎT�;�ĩ�(������)���A�^�HD2�18D1�/���P��z�x���zY���r�:�I��",	���a�tsW�f�U����J��1J
�+G����� �8P��&y�Ě�ъ>vk}$�G��#p*�̷�Aj���vr�ű�p&��z�2 ���L����q[A��m�zO�2���"�[�!�B�4ZZ����+GLu���h����e�uK�&�2$%���S��YN�wJ�y�����LN��|,|h�� '�<��d��HwZ�����.ǖ��y���'>�����hw��<�Y��4�ʣ��Q�P˫��F'\� 4s7��4�o�qK�8���d(y<=�Q����S �A'ix��V~;#l�T|���FY����Q1��Km~?��˖`p4�(�)-,�n�	�v�)�|��Q����'ih�٦���J��[;�I֞�6���>6,��a���D���`g�^&C���*��]m�����w�P�z\^��p3ު�N�'�Sx�������g�d�>�'�W�
��x�����i�5�Kɗbt xb�6Do&q�LgN�����F���ak�nVȾ&��ﻇ���[�h��$��}X8��l��6d7�;�~�e� ���OBXT��zы�2^YF�F������_/[Z�+�|��L��[q�[���+r�I��NX0O�E�螃�7ڸ��(u�	s��[���Ӎ}`[��\.�s���Q�3X�Y4�L{��zEXJ�$��G�hz8ҧ:�zj��m�	Q��vI^�S�a�#4��)1Y�l�p�I��#�嫎�h��JaI�\�<`�"��ڲ[��Y���m�+�nALPQ7 H��o�HY�5s�P���	�fJeu}�tN�`k MDVU��Pqnm�z�"T�TT�@�
���oS���r�N��h�\��@�.>���砞$�¥	�dARK�EA��[=P.4�����@�y������)�-S޳o�RI�L
X��jPx���^73*���<�ϊ�}r;����c.��k��+��<N^���Ը��RF��C;)ES�I���|���׻��:K�,��x' 	39�uP�
�n�Iz}����R�c�$�~#e�mx�-!͎�pe���x��[�@�}l;��BD��[�E&{�HW�G8<L��y�!��R�ՠ�h�>4Ñ'ʒ�L.�I
�;���I��ǚ����Yu,G���r���n������� ;P��ng�d��ཡ��Ig��Ro#"hr^�:�r&'4p�6dG��W�ʯDL��2�J�iS'bg#8�v���[ӊ��F��4�tͨ #~`��{�u�_._�(;����;���@=�����i]Ŧ܇�U_�s ���"a\��8d��Φ}tr?���M)�Ͼݩ+mG޺�%�c���S�:��$ $���2���z�ά�f��+놥dTE�s�m����R�&Ⱳm��!�u)L�2@Ut�4�ZQu?�>I|'�C��fD�`^-�يG9]鬼t��� =����Q����/��7T3wd���6P�TL�|Kjy\�c����Y�y@�UQ�%>�1�%!���|����O-c�)vv�6�f�PN_�T�l���+F�<�_OKʮ���JE�˨�w�����X`Qѭׂ)C{c��m�M���RU����}
�NU���9�$/��B8Y�wM����%�D�=���Z���~F�ß9�*�HxTlW�����2����4�կ��O�����]=(��H����K9Ϥmvm��4�u-Sȵ�bԇ�m�3G�5)7<�g]=��zO�q�� ���d&�+�Z� �B�yN|��^W�53<��6�GJ;�͂����X�y��u���4��H��)x��?mz��xG�%��"q�P������`���>�r,����2�%���/a!�Z�`�p^�^��Q�G����/������V���%� ���O>�Ɩ�NN�Ts�u�ȴ!���ăA�Ɖ+�!~�nkZ�R?�h��H�g|�[���*��-ӿ5.�e.{@o��X5�G�0��3��Q�(ɷ�m�J�J3�7��ѱ�˸�����	h"�4��1�(������/N���y�|�o�*��r�`�F��Bށ`�%����.@i���k
 �bz���� ��u�Ъ 3�l�⽡�H~��d9A�JB��-7�|K����Ĉ���g��l{#�n�`r�u�ǹ�:�:�&�i]ugO��o�2����T<?,/��7���`��Eh�����4G^B~�c����r�zڌcS�jM�hzd��"qYlo5�Az+�����ن��Q	�4�k0�s��ᚶ�[�bR9"*��Cx3/ޕ��S�����p�Ƿj։�J��(����#���><�߈sm�p�Vp���kɬ�n�۰��!�+�̷q��x��-a@p|D��jB �U�7�J���)�>~���F�����G�|@;����ָ�y÷�Y�|���_Γ� ���. �}��QKf���R�k4�����Ϙ���fI�yf@G�0\�j��U!��5���Z̋�D-���'K:�ʽšHZ$L��K;p)2�\6� d3��!6N��@N���`Z((��π"�5�WŪ��t$��� �x�4���j�I��Q�G�a����l�ܔ�뇸��O��Zͬ�M���op�����:�$��:z�-`���"|R���.��g��� +�����Ē{��2�[�r��������
�C�X>�n9����6�Z�ư�
D}y����9ہ�f���E`��5B:���8	��9���D<����x/\
��م�H�a/�q���y���V��a���en���:�ɛe/aQ������#�s�r�7�q��ʄG�E[guX�����<�'��d��Z�Ț��''q8����V�%w\b�tz�c��Ζ��w:N�!X�Mu��'a&j�43����d�8�s�����8yެ�q���8{w�|c�1
�- T�}�����G�8�Ff�b_t��2dve�\����ُ&Xm(��l�<=&/�d��\�g�am_���Q)a�5�Ew�x)3��
�>�h`Bp�z/s��1�|�qt��S�;�d�\��󅌤XD�Ԛk�ߘ��
���%���r�hē�	�c�X0B4f/v�~���hX��~}|��1&���Z��VN��;Y�}'�ؖ0R�"N�S.�-�W0rl�
��F�ݮYC����l7r�,o�:]kD�X�q��n���~��칖Icʼ�aF�q'��U�x�Og"�N�����5�j¹:�Cm̓�|E|�{#���p���o�Д]ƅM��� иڂ��N��Ūת�z9�ل5�Y{�}Ƒ�6�[/�#2�p�z)q=y�ߔ����W=��4irE��.<�s���8���`��?��R9P�=uo�F�Q����<w.��̲8�P��A�� ,K��i�3�@'y;uЪuj@���Ŧ��^ftn�3��v.8���wH;��@�?M�{�L���u=�u=]��|�g���i��m`�Ҹ��Ό���X:��c����5c.n!��t�'tu���&	}z%�8'
\{Ⱥ��͸��R �QŊ���^�
�����r���Z�jG���t*d�w��.u(���M�Z��o.h�{z���%�-rT`Oi�_�%�.��LT\Q��Hm!^��Qz�n�h���V���Ո��؃9�bƮ껳�oc*�>7omǝ�ay��jwG��J���yP�RDtJ�LC��#�I<U��OLi�k<�����R�V�����IV�,���/:����L�T��ƣ�?0��������"�j�?���	�{��|$��apj�t:�Ӿ���p;��<H�4�|�R����4 y��W)��41a�˸�)� Z����%Bz��˅1�l�?b��<�
�cB
�A�j�9Eω�9e;F���l��4�E,�ە�9�}�Ҟ��A_���E|��N�ާ^U���.v�'y�{d����4��P+���ii�A�����ش�)�,�#��T�W�^�7V.C��eCɻӎ����"����]���:t��/�����f~��Q��"�2#���J;	��۫?�:��O�q�����6}�G���.��B�T(+�:���R@V����%.�iv����K�ƃ]�ku�s�ޞǻ�7i��u��'�;?���,�C~�}�Z,Yԕ52'���i]4��(Y�婿Ua�LU��B���@j���g��p��<>P�>�D�1�0���|y�:�^�}��{{��ȭΔ���=�9��趍]�s ���*�=Y��@)��U=��CvY�6%+���U���qa�+����q�|���*���gl�lKnT
8|ɕ�����RG���F�>W�Uy�A�Xw���z�h�����ƀ�(=K�;�^iI�S)�#���$�4;�G�/��&x�%'߈I���*�:q��`�ˤ^o~����wo'{s�8Nbq�r��3Q^)߼��,��t�7E:Э��@���I�e�I�x�.lQ��!��2a���D[H�!8��f�#�F$$/EX�?h"�"��fԟ7�޷��)������{.��ws�^x�r�\������
��{h�-n�h�{i�Sr����mmi��H�[���뫬�`��R��:��������S&  ���[.\<r�"����1���7�����j����q9���<��[�%�c
�^򄱃�Jl2/�J28�SN~����|��a0�6N夶�q'�J������!C.�
��e�w����,n��O����D���Z�1����v��ĴÍ3FA��ǋ��^����p-����3��ܪ�m��d�����R��������s��i{z7���y3a�,��R��#*"o7V�������T᧽n�o���g�HC�>��NɁ��g��Υ���6A�Q?�g��V���/2��`�K���D�bm�0�?�ۭ�����b�{z����x��'�K�����-����&P�l����N��i��#�	y�T�a��V�� o��&���b�W�q�\�%K �CR ���a{�P3�Il
� �۟n��j��mY�o�F�e�ex:(9ni$�Er9�}ƚbh����W��~�����Kd����<Eg%6��),�ۂ�{�y*�8\
�T!X����ט�.|U(�{�znG��wI|>��sb��pՂ\e�z��&y���Aq&ע�0;��!ל"��\�Y~�:ngF�q�byi)7׺�2�Y0����Ȁ���׵�0��iCc��Z��N���@x����e5�y�,c����6��X@;��R�)�e�z����N�ro+x̏�d0������d)�gC���:��Y�|�pK�+v,o#|h�"Z�<Jy�u/���*�� kV�(�ġ$�I����o�[���n�sΌ��l���ä�t��JF7���W_��S˨�=���
�0�~��BB7|������ټ)y%d 2�[=�@h����g�����_U���f��u7����c��"��)�V\7����)g��Mu�%���U�[�@a{^��z�y��M�[庑�O�^��f��S�TK�$ɚ��mQ��D�O/y�J��00�"������p�y�|���q��g�b�m�t�u��q+�ԙJ�*C3�d�����OL��͏�S����L�6%�D��,}���U���z�`!�H3v,m�==}�,_or=.�C��<g�)b�\���\Oά���1�5�`����	��c��HW5=y�����7�(�Vj��i��B��'t�f�W�����rݲJst"!�z�h�J4;��C�6t��+�.�!�c�^ �Q���e��8�%�震����PB�L�{H黰j��tf:�/��H�m��~9�
�/��iϰ~���|��ӕ
O2���7��ˍZw�%��0��ќ�D���[u.):���&Y�u$_�V�ŉ@��$e�#����
cx�p�͒x_@�v��g;"4�,�?<�5.����:8: 3L$��+�n���x�c;+&�.��ST?m��z'��k�u$�2E���+�!�z���)(*�I�$,v�L7��pi�'�wyӲ�鼧ܲ��
�n�a��l8;U2�$���PT���uk\�;����,z����Z1z)�D�>��1è�u,*{����Hoz�k1�
jn�D+��{��M��4h����&�[WN ��qm�x���d�(�TB�W�)�2�>��竜l����(>�5&ǀ�y�$u,�׬ʷ�ؚ�����Of�c�H��,rf�;~��8#K^R��	�)�b�r�f����YƲ��R�0�jd����M���I�av�(��=���2m�悄@����>�[�Ύ.�8%ԗu]��أ�*:6�.zQEH�
:�K���u�7}>����+ ��N���:�����k�< [�;<�1��m� �(���Yҍ�b�"�>��p�/� ꉝ��f�1�G�,�� *�IݜA���%E:�f�CN��!��v��I�Zh�ȯ���C�gR���b�Bհ)|Y37�a��ޘ�����ȟC&P��a�[L_�*	Q0�u>�^�t��S9�d ?��l�����V�͹��ʞN��̦�9�JV�����5���J��n��ތ ��4V��	�mC�B�Il��N����gW����R���� ���������0�Z�VbkP\�g^&�l��[��B�:S˘����L���[���g��֝¦9	@�F0�w4̚k�q6������?�E�r7!�c$���DZ�B��.N�T['��9E�K�㤩���2�h5��/���=�����Ǻ�s��j�k#G@_/�Mޘ��Լ�F��]�����cv�2�4Y�D)FC��"jS���Ͷ>I�4{�Jg+!�y�(�r�@��t]0�ј��fn�Mtl��ǩ��T�U�rB�u��K�F1��݆��<�������6��+.�(m_������T��n �Q��ǁոy�^�X�����q�U$���]�K{�0���9T���˰h�T��IB��Z�(IYJn�9M�,k��7��P��Š������K�qI��Jf��{7-S�>j�K�N%�B�33H��_"�u����˲��ԛ~�I��uxv��Q� <�Nn���۲��Tn�0�֘\����uY*��a���K��+O�Y��[F���y���6Ǣ|��L�+�mص��_������)֘�ǆ?CQ��8�y�g�w�}�֔2&��8ƫح�
.�y�5Z4~����Aޠ��e&K�m-����ԣx+���5&z2� 2h�n7�.ƌ\���ݲ������C�G3�lP�{���T�?�B���SIڦ�~�4�~��9M����B̥�R=7xD�9*��7V�/���\��㛖�n1���]I�I>L��jwǋ�P��`q{�[�R�0*���X��1����e)DK9����.�g�[�N�
�m- @��<b�hoq���~�H0C��Z�  w�		��I�)vn���v��>��Xr�a
���oo�i�,�9!u6�����38�T� .ho��.%��G1�B�:�y$A�'�x�{2��^F1�=��}9,Ī9��~:J����3ܭ,�[��=t,�U�=�Ҙ�G�n�%��u���9+�M�Y���{��ɴ9����������ғYb���K��.��_#փ��8�?�ɒ-kǭEd$��f�t`����^��mFZv��m"���(I��e&ց'$�`{ ���{H�n��st�^n�[�C��{�M~�[�H�"fq�	|�F졿�&���AȠy�|�A�Jϴ�!_���&:�22���#�,�7� ���a����0_��u��,�ֲ���iv�(�\�{�W�.S�<��zl=X~j����ƨՅ�ᅔ}Z�~�*YЅL�i�<�[M2⚞�T�լ�����М��� &����V�;�`lL{�W}E�;�R�Y܀�����z.&��z�V!{w̮�b��q\O�:��]��
�YVۦ�����"��( o�xh�v'�&�����LB�Z̈MLS�c!���6;��n��#�X,�7�Ig�d�vǶ4<��5���a�"p�V�/��?�I^m����؍��p�
x�G�)-s��1=��$s@���&�E˰5}��6��;�þb�` X,k�����;�5�&���s�m�~���9�p�A:M�`��\3�< �'��R�$Ѧ�����V���j\!�9�u1�E-��o��p���C �*��I}�SQ�F��0s�9�j�\y�}�b=�!B�AS3�{x�*5��J8TA�.�e��bߺ�-Ur��C�K�3�^���q�x�5���۷�f��8��[���?���j��Y��!$x+�����WƋ��zSEfnK��M��:����[2b�wW�V��!Z��Ei�]<0��2V^�O���X��B۾˩�)xX
1n����e�"҇^�T=�N��u��]Λ��e������D�\=�h)� x@4uz��6�M ��f��f�hGƔ�h7�վ�ڸ���u�钓�*�g�_V���IV��;�,�'�%�+�a�����oJ��Py8$��C}��O��@�Z]�R�n��br�K}k[���ڍ��@�>*uǬ~����<�R�U�k֐,S M&�x�V��x�62Lxm@��W�N]>G�+tԞ��K�}�[	��(�����O,v`9W��"��֢�H��o�%�#B'*�82#:��w�� C�)4�E@�5�
^��jc�nhzC���8^%;��rˤ�(���sb<�.��6���_������e�Rx֭�=ɟ��(a��+��l�t��[��^<�4-�`�w\���O�Yx�8�5��+�F\/F�T�W瀿�;��1���@�ٜ*d�z-���ä�]*��ˑd<<��Il�ꓜj,�zNɅf+�$��;���dAdڬOe��^����+'���|W���opdQQ�15�8�6����c�ݘj�7�y��s���A����H�+���ˆc��S�,Z�p�Lg�����fMQ��)QX�}B&rE����v[�a�\1�����=�"��b2|�JKŏ��Bp��6�7����Cn<L. �̚'�ݘ��8��:j�[!�PA|�덆&{�$���[�5q�y��4%��O��E��)��|6r4f��*�³��&��H����Ʌ��iE��d����U7M�g3�N���M�
R@�4e*�K1���=�6Q϶p�4	$�����\��^�q94Ql�5�ՠ��f�ty�ŁԀ����ݻ^IH�_��X�h�f�0!����ގ�I@��v\'%�FNIJv��>0�
8��m��K��G��r�З_�>s�e�H���Q"St2Ͽ8\��i��F��:޳t	�%XB��[^����m�$(�E�	�ωMe�P�쿘�S�P��ܗr����79+���^����>�7a�ڥ�Fqi���r�qP�8�)Ĭ���Q�eh8�Y�����g���7�o��Uof2�V��/J�q��e�p�ZLr��A&�e���(�Q5W�E�<���i`��(��2�HV�C�*�n�WMi��|��#=��l�Q=�3���B-�/�
O	E�}����1Q�����M���v�d���	�J����ht/p�Ct,��f�@'���Ӧ|�
N�97ﭣ�G,�Eu9�������������VX�#��I�l/��}���0���4�I��+dx�T��[[̨�V>D���N�9��?��.�,'��g2�O)o�
��%\�7������tL�l���9(¦�9GR��c����I�n�(AM�GV ��0��ڗ�q)�ZGϪL�Q�ǣ�V��Y[Qg�"�_������t�3�9����~H�x!�<	�_�k, M&��H�(y^$p{ˡ;����]P���ݮ����T�a��s�����rӅ��Ds�̎�ϳxIP#�2e�\���B)�Lݓv� ��F@��Pz|�Ď�Ϭ��c�0�ԩ҉ ��|H�B�n:��CO�y�i�� �?�0B�tA��y�>V
��4��������n�%�W-�z���:����^��:1v��h�e_���_�h$�Kn�_�O{
�������t�,��Ҋ��޿�s���L_8ؾ����S}B#{RHaJ|�_^���Q!ax�4�O�-�ӤS�75���`�*p@ۤ���
rL��I�xv&�N�Պ�2����ME#�a�=���g	/�o���(,|�{���Ъ��@�R8����#�H|}^�Z�2l�>��A��ù� C��D*5]�,�g�@���j2���@縸sc�=�K�F����B�B�� ��~6+@m�i�ѷ�1��b�i���{D8y�wd�(q:}%Cb��孭�]��E^���Zq{dS��j�@�m�!�`��x?��h�\B��\�J�{�jk�m�]]K�LvB���'f����c/��PCc������Z:����r��8۫��Cٻkq�u]-���z5u8���C����OWg�ֳ��;�k��̤ˌ�V�
qX`9K�V�w+�qL{���{��X�H��"�Z�$*4�x@=Bi:����nFP���c]Sy��GG�5My=��7uf����KZ�͕l�� �Eb���e������̈́�T=^͌N�/>�f��>Vc�2d���c^u](	�R�G�k7
Nu*҆��-,?B���_+u�\�̕����IW�h3�K�}�eG�u�c�+��E���.5}���6߀T�T���"�[q���*��[����T�]������m�@�P���M�mv�ӟR�ʒ����o�lwd�_�in��Y�1���Ѡ��u���Y�n�08���Os�r���=<�b�>#�ݐ��tB����A%Ԑhs���JɃB6�:�S%k8��-�c��Ⅱf�g�������l|�� �0.�RZ����=�_̵��𮶦�c�h���*�wXE	˹�GpMJ/�+�Ќ9G�����cF{q��lנ[�Z0��l�E	B�R�V��"ANE7Өىb��0�-a�O��rh���5㎖�]ۙ�axMw�A�4�8h���#�.��Q��1�!.�Ai��R1R�ق��|�]	��� y9�mgy�Ml��T�N�f�
�<�~�t��34��������0�*{�q�aP4�$}�+�4]r߀?߆��i�\��.'Y:�����ZM!��p�� ��؏�^��2��Gi�h����i��]ps�����q@4ߺeL��6��Rm+kEp2cn�W�;��ni��(@2����s��,Z�-��@�uv,a�t�ի�^��2D���b~LZ������R�R�Z�ӏL�>�v�����PǤ�j��nQ�(�����*���aѭ`(���&��m� ��x�KIj�*��� �u�������v��]�ʲ�K��J�A��� W�a7��O|^�ԣ���m�ILɯy��k[��Yퟶec���u��K�>|D�<��W(�Q'!��D�>��9%���:ylL/�#��d�ZyC-�2o&��N�k�f�X�Ԩq�X[�-<�rr��J�4�'�Z��3�`w��/�;�)�ZCi�^��Пy��YA=P�K�]�	3@0n����	%'�_��,)G+á���@�%���_�YV�q����%Z��.�i|ϒ�T��G���|���K�3��@^5����z3N7�E���s�[R�Х����kl<k����qe�0�蹃ʜȼr��f`��	�����FX�f;V)��)@3�;I�"7aL��W9N��^"�f�Y�<BI��Y����;򟳊����iLEQ�Ǡ��g�x�F��%��HއO���Rg�����9�2��OEv�÷\M�|i2����'5_��t$�j]�Fk����m�3l���rM�`�9+12�wG�u�}��h�|���A��T.<����|[I�_�}z���(��P����g���Y����"p���A��� ����dɴ$9��&��^k(��3��H�ν�k��y���v�[�O��5t|W���Q{	����Y�rp�w���p��;�{7sm���%C��ف7Wt냾�D!��mr�kbq�FMA�����ױtg�ο�bR�k?%�]���t3�G� ��Ʊ���֢'a��!#�	<f��C55�F�yB�;4,F>�_��]E�'�鉿�Y��%m�~/���4R�	u��Q�C��մ]���Z3�l��Xw�מ��C�X�͙D��ps�66�+�0�٦>zKQW$- ��-�21um`�C�DDTv7\���^�I�I��xdm�5��wo�'(]���֫-`�z]��fO���L��.��b�+u��L���wg9���n�w`����}�zG�aAD�����pM	��S�	�5	�{�(�<)U>�ƹrkR�7�?݊3���&����oj@@��-�|j,�B2E�Ӱ�L���F���x٬�hƮ۔q����I�jKiز>xL��l�Δ/�60O�ʤ�h�U���[�s�� hr7v	$�bWj>�&�4�=��������x��Wm�y���[�Z�ϸ\�$��������̋������T8j�T��:O�Y���x�*�rO.6�V
v=P�2t%ʧ����۴���\}D9��O	ʺ�s{1,�[ɋ�ab��#y�W�!_�5��s�	�����=���^dcIl�����XoQ�Ǖ�hqa��[�S��(�R�1���Ò���/��@k�Wp'�Z(��n���C��a\n6U�k��+��[����c`�]�3�T?:faԹ�9!�v~.`Z�.��G�8U�`'�+��i�����<��8��n���}۞�p�Ƣ?~?�G���a|K[���T ��7�D��`��	�KzЯ��B�wr�c����'���i���bO�Q�>/+���~�n�ɼ`ɩα�J��K񁟍����Y�ZV*~l6+�a],�Ɉ�I>�nI��ѓ?(���G�;l��T$�U�o�^����I�d����'�P��@]4nP��Q�k�Zxi��B�[b�E�>�6鿧�W=������xl���޶�]��Ў�WG��}���-�s����:F�1s䱴���7�*�ZdO�S~�P�α5��pɼ���S&\��]�_*�M|�e�P[p[��_EΏQU(v��q���)3�>B�����d8!�z���dݘ��d��X��o�1��P~�
5���E�8�|S�mz�~�3��T�Xm��U�A��z�H�<�����cCT����qo�³���f�F�A�kv���j��$+�p�2ZQ����M.F7�}�,�r��]�'vn|���sſ.J��p��?mҽHQ��ɋ�Ywz�u>��@�=S�p:U$������F(���3`JF58M����z������k4 ��]��H$ã�q��`�"a�I�����O?q�+&�`Kc���5�,P��\I�ZYe(�4�Q�H��Ö|f�?����(�b�c�꼤���a_���k��w�l?K�`ZC��eo�q
��0��������=�$Η �q���f��^b�Z�˰V�K�i������0؜V 4y�")�U0)�Lj:e?�^����o�֍�F��l��ȫWR�c"pJ��Ts8#V��(	�-C�EV���l�60����Pi?HQ	v6���PS_�U<z��2��@þ�oי��������Qr
��}CkR��[.Kp���⯔"X>�X�pYLѩ%���KΕz��}o�hٿ��i D������]f�2,ez�����y���Q���N`N��[�����N�a���K��*�׶)��t��뺤�~��%V��	���M=���9N� |jb�X��.3�J�J �/��i�E�h��=��^�N����d�$�e9���7<VO%������eY[B�E����Q�i�F��8S��9�fkh��9û!M��T�X�h�~��ÌBڳz��O}�1i,���3?C��k�n]�F	J>ʤ`}p�%���O�:x�~��* ?̣t@����=�<O+hr撠Z�N96�4ݚH�&���#EW����X��
�-�:*Z[_>�k�����Bب�{*�1�Y���`���益�&@�n�M�l��
�pV	JH�s�����T+��[Rut�^?.�O�
����"�"�t�P���?�l~�?׾�k�G(L5~�a�������V�����[d� ,R"6�H��Dk�l=E��#��.NP0~}R�f�UȺb����U*�9�x �#�C�i�[7=�g0HԟX��s��KC��	�xL��2Q��5k�m�OK���~\�vZ�~�#�b$�A�y��b]{��[%�� <T�1����b"�n���sJH�J&��wiW�L:�GA�@�*�bg푶�� mZ����mnDe�W�A��}>�Bz����̈��_= P� �g�)�c�÷V��Q����|v��^�'1�DZKA��B&�G���_VKV ������] gT���SmhVE��C�>��d�`�A�#B�כ��@�=`�FD72{D��9���7F�`{�ڑ��#��c�X|�f]V>�ӆ���gw�{㺷��P;�H]��(���;���}+ܐ��/�G��?�������. (�d
-F��������H{T)�n�@��nj3RW��y��������E��U�͎���oj3��|M�Z
�z���h�E�6�}���*��v�U�%3�@g���f-���<���l�1�;�=��Jp�S�H7t��������#[7b���4CBiPg#D��ɚI�G���4q�艖�[Ey�b�U���l3,�aq��c�Wf~�ơ�)�Hľ�kl��% },�C���{�|���%z'B�]�4��\�%���e��QA��nB�<%0c»i%i����1�`�gHi�V����q�A��/���?�1i{>�9O>�ɾ$� �̲S���V��N��OHG��M\^�kn�25�!�n���&�#E"��x��b��'Zc�NlU�8	2v�+���|,��%��_�NV�t;��Ŏ�"?:1��'��7u:��Gp�D��ʝ˪gCo�oIY�����_�������«h;����nD�[�����
S�v�zS_)���5�c'8��w�ҍ���p�: ���:�bK{���\�njt\�G�c����=�v�쒪����))eq��Z��M�P�<�^9{c�Z$Ng.џ(@$� ZU��e2qm�L���!rx*R�P�q�L9u��6M#�R�LtgV�rl�3�l�@�!��%�z�"�ƝP�-���F����:���	���ʲ=)a$�#^�.�#��b ��]^�$N��	�ϖ: 6��gSy�7�&H�[ 9ɾ�E�a����bX�5����Uʅ��3kz�"�dLY3S����tڪ?��^�U>	���C�=�&��;�K'EeX��Yg������d@�^,/)E�t&�?�D��Q I�����l>�O�bx81ܳ���@j�Aɘpj��gދs!71�H�U<���n	V~P���@?ژn�j��y\_/�X�2�M3�1�1r��/���F��d�W:���طu���N?ږToϝ��G�f�.�C�id*CSM���W;�DoPV���a��|2JMr7����wpq����&!U���ϥb�ӡ����j;��g\`MX.ct�G�wP(����u�|�ׁU^U ��ܸ��++pI�U��l)�H%�H�Z�ֈy�"�RV��/aN����<n���]:=A��������y�qJ]| W�˨R��\8�f����c_St�C,��
{�K(R�4��X�@��ôD}y�`ծ�n�H:Il��>U���=R�{(�B�Rsx\L��W�<�����:�^C�N����zFgs%i$u	�w3�I��A`N�E\A�㈤�cTߙ@<@1S����9X,�$_5*�,_}ȿ��'4����!x��R�AG������  �O�O�31�W04�B�w2$�&�qU�a]��4�]��I���F��ٷ6��	UTU�D�@[L�<H������]Y>� OJ=T�`<g�m�;ׄ�]�>,�4��"��r����^�l�05]��F�oMJ�Cts�:������Ox�b40'U3���Z��t`7��p����G JG�K�����.bOd�"6Z�� Y��W�=\Ȝ� ��6�vٚl������/尶���˟5N��r%B��7�}��?p2¡O�:�H7%����E�b�BcQI�`h~�����$��}�����8�,{s_f��d(�-�������÷�+�hw�V�F<�n��
�w<鋙�m�i^��()R� ���F6�1_�l*bFͅ@��3���7�� �&i��[�C�S��B��
5�22�f+�q����AC�����-������O�;eC�Q(ÅV����ި�ЂY��N�ԩţ����%�<����d��TL�0��+�������0�c�f�0���Es��H�f@�M՗����s_��L��
v����-�|	%5$��7U�l��;G��i�GU(�`���"o�'7+g(C��	�zj"Р��s�N�c�*�~\��'L��mo�߱��/	
r��8�>�^���N�r�x��}ۓ^hd���=�Ua��X����+>%W ��'����pC�oh��8���
_;|&��^���?�;�N�U�44��c����oY=ע�ݛF���?�jv�
O�YPV����ƣA2S�.�x�k�'��4N��½H��e:H�&E��ul�V�H������G��Ϫ�Ok�f��߻�C���s���p��/sR�iByx�x&��S�9`�["�!�!��Pz�R=��-�};�p��,7�u�1&>"\�L_�Ն">b\bO�B��Y)��=Uȣ'���֧��%@�o�B�S�JLCz^�ߍ�`��b:�tN2� �5�lE�8��e���6��Ov�֪�u�w���B�6��ą#\#*�3x�P��}�{8�q�d��0^�g ��CX�,�yd �l�b$�:h�m��ʏ�m	9e-��3�����q1l"������ߊ�P��j(}�ʗ�E��X���G���<�ʖ�����ymz�t~�
���)$��I��p���nQ�\2�lQ3X�3�.5��D\�n6G��B6Wh2�y]t:1�y��I�""�/K���� ;���SWR���E���>�;.kR��,�Q�*�~���Z&"�����zI��C�s����}	o0��&,�*�zɆr��l�J�=�|Ʊ�S*�ڭi�
�������G�N�2o��,L��$�9�w]�:;T	�����mT���F��:m����vEt���������2u@|���o������9/� �2��6p���N�6B.�����zݦ��w��l��h���U4��`,~�PUd&t��^G�x��_.w�R�IQh��l�v_*4���D�M94y��K4&<.�V�~!ވ��<�xr�͒�U�ΊJX"�*���� �.�8I�}�(���Յ������}������W"O\E\�pM���ܮ�Xva<Ծ.�xT/%�-�����u�IZn� v��I��{���� Dg��U_b�y�6H�f�.���T�bv�/ �_���"+Io�����y~���Rv��;���u���~PQ%�5��g	y9*���4���0����JJt��w���NiB�A�=����z/y�b�~s@�l�2�N7�q��_�&s� �8�\�V�U�2�%!���o�iԸ���F�T����ŽV��`�ʅ�~1��%��<q�*���L�P8"�Te�+m�E�]�GG�d�%�:Į� �w̶f1�̸�aԶ��i0�`/T�cj�52��Ҋv�U��_�RӞ�tf/�jy�'��Mώg�M� �͢�c����6 M]���W@
���$�d���h�*��M��1?=����m���B���u"�`�V�7�hh�}y,� �����O�jfJz7�Vde�R��.��\���IQ�|�A;�_��,MX��*�;�\��A�������)ߠ5b$���D��Gd�cfW� ������V���B�qF��'� �.�� m��n��7r����K��S��C>:�r��A���3�����=����d��zzj�g�7&���ߧ󎤅^]��ZSG�A��(.�� ����uc�بwB���j��V/�]��š^��5vV�fyas�D�&5ܴ"�bJ�� LЋJ��2,OI%ޞ�)+X����C>�
�x6]u�L�^=Dl�>M��7A�Q|a9[g�a�.�{�t V��+�����Q��r9%#c��:ǜ�܌;na����������Ep�z#�9�݉�6�l&���%p�dat��h�Db~U���gc)C�{4��䯱n���p�� �H���3��y:��Rk�+�T��dkKx1%"~�
L"1,P�-�o�V��Ⱦ�ĩ�I���S;���l�4ȏ����e�*�G��E"����r=�ϔB(��o[����,�/���� ���!䳶M�W�s�5,a���	+��:υ�#����HYe���aIdI/�X*�$ d
ҥ���p�)�т���_eU9�M�[4�3�+W�`Y��l�re7p@�n/�}�(9�6p�)���7&?��a}���iIϕ��āqG�����^�(����C`�/��'���\oJ`�u��қ�1���}�-���E��9�v�r�+$Q��O*�Dsi�;kYH
�Em"����T+~��y�B�ݭ�˯E$��P��~�2%�dUk�QZ����_0B��#��_նN@N�{C��c&8*@����`�s$c�
BB��cW��C�����)�:���4��W��#`Ci2��răy#���rZh�3=��#�=B%���J�~V�/��a#�{G���� [d��n��8��&�Pњ�U�
���Yu���Tπ�Vm�oC.���cy�,�y�p����^'�M�Z��[i�ZY-�t/ʘBP �b�0��:s���2�̠&9uY]�
H�[��J}�T���x�]I�	,�5�T �m�̯�
D�<�~�l�#� h�tE�eU��l�w�:=L�&ŭ�%�Q��"+<{ķ�5�UH_��&������ �9���;��E�� ��߾���SB������$�V�/�{WbIB!0��/�bY�lzd6�ī�X��1EBH/)?�4��\��ɖ��	���+�t��w�3�RW5��h�2L;" �Y���=q�����Z+FO��ɡ�Z���b�K
�q�_���$.�L�ƙ?"�R�5�?�0���?`2]i RR�T
�Bc�r�)>�B��>��H)�`�.K����S���78Z�/�����,a|J�u�FHᑖ.�a��\4���؈�
�5���Hx�>�7&c=e4�`&5u'ٽ�[����A�k�`c�XDpK���	F�`ә���aW�v���@t��VO��aWhY�7~�%��M2Q��}F��,�	ǡq�>*�1$}=!��ORh�+�5S���8�]2i�:�̏�*�ՋY��=W<5��M�y@JQU��;r���z�7H"g��xz:$� ��h�|S�����32���)@�r7e}}�m���5�;��͟L���0OݭA�F��WaX��1�����P����M��Vm{�CJ�P�+I�ub>�=a$4��D��$���v�W��O�q��m�d���y��/���s�0����:�[q��ћ�إL
~oN5� ̨I�i��8�+\|"�qY���dE>��Y�Q<�K�\���E�%!��:܅ {��U1v���7�=�rX���:�fЊ�enV��Q�*FϏ���ɡ��EDV���>9��%�(c��R.u\�1S�]�DG������.�OV6�4����nwNB��/�2��u@�@��Y3��(���n��΢��c�^&���J�T$�j|^�+�V�nU�#}S�Ɏ��ڑl���W"Ihx�B���W#�5|�vbS�آ~A���4�O�Y��K��0��^�����|�&cx�8@��#d�Sb�F��u�k�U!�m"�����Vrn7�(�tDZ:�VS��`�-�n
����s\�[��ɸ�<�vW{<e�(���3Sfr7-�--jJ鉎
$�"�3ԇy�b#��?��5\����P����<t	��'W�\e���=� ���5��/�h�v�ׂ��|W�2�L����h��fuC��)Z��ƭ�d�ϵZO��7_ ��}%ęDn~�fE�]�1�=�[vɛ-���q�
�s/��D�A�v	�(�0<�`�0C����+ F;qmM����p���}c���[x]eA�av���=Lnd�i���d�c9Ͱm(f�?뱵�w���e�(99�a?MA��N�� V���ţY�-��k�6'Tj+x�l�Do�7�f6W�V����Lt������vc���\f+�i��r�+�Ύ��N+hs(���ef�?[c.���]��w���#bM�z���f�n:�C7S�J6��7袖��dU?t ^��C��a��uÙz��Π���A��5Ҹ�je2�Tm�� �yP�ar���g��������	$�_n�G �������z��á��07����&�G�*�]SMw��
����pۜ&���� y&2cBQ�T%֐���/�1wZ>*{%9��a��Pp�B�Fd� �B�J#�9��:*��^j�Z^��꒩E9.��N.��)�Vg"�x�œ3�
�I���0G�0�<�1
3�[�� S�0kG	�Ml�K�%��������U��R��B<�DC e���?U��pcX#���u$��H�W�I���k���sRC'}�������F���Z��X$�歹B��C�<�!���c=��.-�6�lR>�|:�f?�Jh9t�̆�IN�=s�\��8)FR�?��/��={�Swo'tY�ך����s����)>5�h��\���ӑ��
�/o���vX�OnMH�rba�r�Q��xI��]�<`�%N���>���p�Fpo���z>!3�L��)qi��vQW�.\���
�<,��A����V���2p�Cql�6�a�P��������m�#ְ��Օ='܏&�C
!��������Iw�Ȏ��4��*���I�d��T�{�͑8D{��\.��/S�y��r�^g�k[ܕ��#p'�o+�~���E��(ˑM*�����A��.~9�'�w�fO��űp���|'�L��-|�L�š��1Q�9�#VW�Pu�>��m-?���ÿ��p�Gק�h�s)�>�9�M��."[1�C��nJGwyd,��L�9b6��7k6���=D�A*���Q�$tPܚ���}���i\�2��&���.=RFvD���B�N|�壷=��yW���L��&��bmXKn(�x�f�2�3�x"����k͏W���b@��'2�E9T�v���]C�,l���!w�U7��:��p����T�/`.e���a�c&@�C�|s���!�c�)O�S�,{k>\#��yl=�>EnjoI$�[/A�a�h=�QJ'������Q�xc	F��\9��f��>ޕV���]ﴘ��X��[b0?���*M�O�'�f^��/J'N��wt���R����%�b/Op=�i�x�W5���e��Bg�f���2n�%�/�*��:W0Ѓ��e[�����
�l����>�!�U��TJ�;Y>`m�6V��S�{+H�B��G��yO�I~yh��sϸ�8`T8��z�e��M�<��4?pFY-R�0��f�}"�W�2��p�Y����zXV���kSuZT���$�aӤY
��P@�*%�`OP�1ؘ��	�:^���'V}`�
����0�m��;���<�+���y��Ev5�O�[)��iQ����M�g���\Ĕ���B�G+�T�- ԉ]e��'�ѡ��{1�:6����K&(Be��G�Y�D:��� ��!˓3�Ո��D��h!��Z<�Sa�:�y	��9�j�:y� N�b.���	~_!��ѠH�><M�s�(7�\��e�V�����
�"N�����!�������d_lA�US��͚G��][���2gs�>3_*!�m� �~_��/����j�r���͚�I�?یg���������V=u��w����j툒��Z��r���iO�-��fT�j9�L���X��NF��iR��*ʶ�ۆF`��n:Y�ģl﫧a!�C;3����$i�й��PC��o�ӻ6ǚ�'H�ؘ0���ӝh�m����Ġy���0x�O���9�ƃU�p�DǾ�$��c:�JRMe3z�8�X/7�����U�f�D��sϲ|�6�#�da��l��z���ΐy-AhM����ѧ�pQ�]M��k����\f�,U��i�<�����k�Տ��<9R��d�2L�p�J��{#V�70���q�]�'��N����j���  Ŗ�u��P�6M<�����9���6�^�����KjX��j)���kQ�2�%�q��w�#�_(��:\kYU��ݮlϭ2��<	�biPN�\��3<���>��w^�3j?]��偤O/o�D+b���@�>Oe����� Ě���{Am�t�F4��Le��U��9����\�V ^ ih���/TD紹s�xi�b�l�l#�w������'��)��F֭y��Ǥr��*~$kQ�a�%9�'�ִ,�'�$�}�~�ɲ��V�upY=�<\��V�H���v���nZ�Bc�8�M �L���Zq��ɧyO)�vQfq��~	Pj6v��tZVG�N$�M8�yͭ�D�tO �k���d����(��Z������'�lN&о�Ш��;n��4j�l@�?��(��fK�`.o��Ay���ҩ�[�q_�iĮ���? c�����j�T�B:�fdD=%��e%Ed�V,��1T�@��S[{%~Ӑ�䅣
��\g�����^�ļ�������\���Y��zA,4��Q���<���}`�1��]�v�ޢs��z���>�R̓��d[���e�A7 ��#K�BpEA_D��x��Vvp�b]���w<��3~ݓ>��ܨ/E����z^��(V�  ���D9P;��g+��@�f#A���p���^�"��v!��+>�'�C�t��5���{�xH	Mb+��g��օ%c��O�t�1[VP^�>�
���*e��c�1{9��W�h=��
��F�!�J81JRp��a�2�X���F���m��cQ	�Z������+��#�!�P�R� �`"��7�5��[;I;�8�6��*<&�h�	���s`��%��_*RU�P˟���y{!lDL����Op���k�����^_�#�̀�M^�����]�0�[f��jJ-�/&1�B����FIig�3�ӍbKR}�l�tg��Jڌ���5^�t�[M&�1��>ػ��E��d�3V�x���b��[�ҿ�^���↋?Υ�g!	�mB+w�����wޏ�%@�N��gտ�gUt|٧^/���I��\�u�G���g�,��)_wTyyN|�:G��������-�	:�nX�t�Z�/�s�X]wlhw�Isz����&�!�f�YN����窳��C�5)�2�g���k�n\��i�I���3�Z�.i��h8�����uD
��7uO�w7��
i����=7w���^�2�U}�$����'�29�R��kX�Gy��b͒���[��ģ<��iW��/�a�}3<d�2�	F,�G����M�9x����B.b��v����U���
'H����2�P��T�dJԄ���}�T��E��w�{(�ʫF��+(���i:P^��=�=_/���p� '�q���:E�h�͟l|�k��������8��E�4Z��0�t<�""���"�	�6V�0�h�_�~�Z�QY�"o�k�g̙��H���}�0;���x.�g�O+x���D��Q��^�;����U�8VUM��v��2quf��>�?�js�w����wt9ѣ�'�0|���G� �4�R������`�"��pm���,��G�M������|�'Q�%�@I��%k����eh$S��[�i �I=c�E{q[�L���~d�՜|�7%_H����{ ���܇a�^�&v�ܾ*F]����snN���J��ꉬWn7�}E�b]|&!�s�Uc'� )�z��\n���ז� 
a�"���|�a*����_*s`v���R�CX���5��<h2cŻ�k�w�"ėJ�n�K�[	��]j����� 2���m�۠�XV�P�'��\9�s�T4v:`�Q~�!v�&��=d����q��p��Tl�S��gv:��ƪU$����g1��S�[��g�MgL>Ǝ�1Go�R������k%H��[�H��
��Y�S5��oN��9y�j"�J)�놵�J�&������Ȍ���a��(yL���}v�f���.�P�E^o��1�G�DM����AD�5�Z�V��h}SrOx�KF�#�[�6ǮR���j ���f�h��z���[��%��u6�44<h�I"дlGr���-�|�q���VKZPi|�F�<~�?����]�#�l#N���i�SͿ��v�. �Q^]�	7{{�� �_"y�q�A���&���G�$�5����N�ْʭ����-�}�4�MH���״p���6)�i��Ά�1��%�4=XDo�o�X��)Qj��h ���8�w:����Ʈf��@ٿ�N�Ghn����x�={X�������S�:�D(����=�)��������g�PUNU��dd	��{Z嚵�/d�瀍�:if�oL���U��<	rp`��K��y[��>�3h�m�)6����f�~�ZU��O����)�c���iU���݌��j��Y���^s��j-ܦ:�&�[��u�w�I�\�Ⱦ/�ۍ]$F���y%U������mQ�y!KOji��k&\�{e��x��;�U[�'��P#�c|�n?o���E�&�麂ʳ5~7�ݣ�|r��}��U�G�r��u�<���,m��t+�������_����M{$l���O�1q/W��q�?/�įф�T�O�	�ZG���A�S/li������\Q�
˿zŝa��E���#w����k��[ȓO�#��^߷����ڀH�E���30�F齣��Y��'����<��?x᠊`M��n�?�e��є����q�*U�|3����#�[�Z�PЀ�V@$I�?Vס������S|o?�P\����n�Tes���r3��c��&�EP�}s�(?/���tյl�"��cк�G�A��OڻnF=)����Z�!�ר��Q�
{@��¶�8݉����brP�%�R���s����REs3A�%1.?ĉ_MOKZ�<D�z~�!.N��/����IP����EӾDPL5� �M0@�@-�8��i2!L7�P��hз�8"ٻ���w��G�h�[�U��W��u��7j	s��t���{����.��c�s
xԘ�W4[�8��-�¯͒�:k�����ҝ���7��Xi��ADjYI�8.�S._����w�K��Z�R��LU��g�㬳��8�n/)/����h^'y�ȡ��k{u�;��v8���x{9��ު���X����vr������5G��� =��q��rd�M�K֢�J�?�t��64�+ &����f=��?��ܪ��ܝ�[�A�%���\&��0t3k����Z;U~'��L7�g�Ǌl.�˫$��p�6�y
,!N�����i��c� A:�\�r(X����ܔf�P$LP�����Ja���p�^��R50��̉nF �"Y{Q��S��u����~[�<���V�
����@�-��J�)I>ڊ��[-��I��}X�@�H5�������܅s��d�J�A��ѐy'Sue��l]*>]��e*#��[@Ǝ�$�>w�����"8Eo����p��c�hxn�����Aq�`%�q�Ě
��ty�OB��'{[��f<c�}|�*�kn�z'*�z���.CN.�ӕ��#�'��)�. ����}��0������R]b�'��d��c>" �2�Y'kد�>����O� �b������=W8�zp3�5��f�0�'� Y� �����dK[�Pn@��P��BQ�<Xx��I�G����ܩ|�������U/�sW'� ]�80��-s������a�# B��ݺ�i/�\����(,>#���˷K>�%ɧ�^^tB?�<H��7���Խ)A��W�o�b�B,E���\}�V]M�Ў��I�����N%?��HK��/,쵿�G���&7����|��׹iM�0w�!���--"d�;�a(@.����A�W�N�3b%Q��X,6�^�z?L~┋�6b*��"�l��1���?�Y4��>�M��A�kkb�G��۬�I�r-b�Q�`eaDν�0s vtz���y�k�P�z�(����nFIs�/IK�w�����/��"��b�I)V\Q�ב�d#t��L�F��A�=�1�Z=qO���cUȥ���XFXy�BG�����1������R��,��(�}pl���b����k��
����j31:!��K"A�enIh/��|}�����%���.#N�����Q���0�?st�#ٵ�|Ĵ�V����s���x�x�����$��5�g/���{t�Zn�
�\�'6��6~X�%���o�.t����@DbŁj� ��6Ӧ�(�*� Cb���}7tU�CR���orh=��"x�����/J\�F�cjwmd�Ȩ7y>a��8�aS�^7x�&y*��_,%d1b�*�|/��n�hhI�,t�����ĳ�"�hx��tq���<�������߸������0K�)B��#���ՏO���ύ�G��O��V �N]g���׀s�Sa�{�9�d{]��uc�Q���n0毖h��SǙ~�A[Df>]SH��&R�Dc)�d��m�������g�4n�$��9"�����<�he�+�(�gQ�*�w��5�$��:q�}�4D����6��-Sxے��h�%�ǤM%�2K�|�i�Ӡ �rwjĺ�&�m�h�_)(N�S:W��!���m:�+:A,}t��������5�8$�~��V��T[�D�[�h]&6UX�3���e�"�������捚� �kt��>a횂x��n��� @z[]�\�:x&V�2�T|�펵 �h������dnb.ʽz�Ir��"_����ݍ��TB�T ��u���N�9������1
���/?��Iq�WٽEJ���(�BP~%iKO����H��_�b�l�{�P�q�\t.I�.�Qu~�� w���Y����,����[`�o��d!싒�;ED��(S����X��%̍�a.7�_���T��>�5n�Q$�����.�nQ���)�����C�+;�����'q$�Ѿz�Xg��X�w�s���k9��I[#	}�����iэ�!~?�7��YC��}Ռ����0>,4^�o�-��r/�DR��P���5+� �o��0$�΁��c����ʿ��n�]��>�^�E�bl=�(���'a��ƈ�pξ{6J��1݃MM�Qk5?���>��6�C��]�E�̵�#�]�����+��s�
Z���̵?����?��F�����Ċ����Ƣ�
С����{5%�H� ]�JR���s�D�E��bC����L��ҙ����Ċ}��o���$�60��0�,>������:�~z�E1�����cC=7a���c�*�P��)p��j�V�9γ"��e k��D-\r������AG*߈8pA ��l7<��՜{�oQ��{�7s��f �ۗőB�����GYJ�~$O�\��]����
�2'(υf������MG�׵8<~���7�D~,��l��@(qp"�Fv��مH�8�'r0'�[�A ޵���"����??R�wǃ	����Ȱ5�Z�ށ�J��nC�YT}��[N���8'b���7y�볅%�����^�E��ԹI�(�_]�i�1pW��K"�!���v��2<V ���{ԙ�|=�������Z�ůK�S�8�3�J��[}�R��-�d�Lj�j���ÊMJ��?�UMb�U��f�i|�ݲ�`�-O��-�F"^�6:�H��qi��T�IU�/u�|�%�Y�ו�K�6�9�]"����2��o�to?r���p�>�t2I7�~#�j� F���ϯ���J"q�5�eY�[r�0]`�}��},����A*��u����&C��B?�@8������?�Y��DlZ��f*F�Z�9�Rh.ׅg�d�N����Z��~��q�;-D*����*;��&EEJgI��z	����'�~=��-��D!�i�C�rF6#o��m�� $ L�!%�Do���?X�]`����M��ːh4p�[���w�카#ȯܴ̼��j����H4�35԰͡�W�n ��)�R?��a=��z��%Ta
~��=w e�����J7�s�@���F���O��j�3�Q���e�Зw�b�_n��~���A%@܌�r��:��xfdq��(6�r�<S�ηt�H�d�c�8Ù��9T���BW�j2��Q"�X�q�V��[4:I�I�"�W	n:p�nd��'C��L�%�n����������(rP���X6��/�0���b��Eÿ����غ�ۤ�0��:��<&�7�^�0P�^��/�����Pnu ����i�쐛��$0�	�ރ�k-�;�fN=�(@
zm>r�����aPҵ����\��7
ޟ�Ts4�`M�g@࡞Ҡ�H�\�{0�)kd�psF�� g�?&~t_+mHh� �_.�'C�QL.�Y~U��{�#dٵ��~��ws"�WA�Q�?S�-gwz4&�Ө��R�:)�C	�sڇD5pq��FR�c�,�N��9h�4�ʖ���qA�*s���������Q �#ً^6���<��(	�1�!���C��Zb���]v!8oeEG��1�Yp�R|������d���6!�m���+���r8$m����1o��PM�Ry�.y?��E�oXZ���
��X��t ��uT�0,`�U<�Ӫ@��;q����8�(=�k�aH|�WUqɨ��6�wA��U��]ex%f��51�U3���ފ��j�d^�R�	��t�Aik!�!������;`���_��F]��"լ�z�㢽l��@lj������2�L`�9����e��џd�� ��p83;
��/Qd9!9:NV>�4t��������>�~� ײz�����_�7I/�]M��z�@�q@R�q�d��k��0��&������ͧ�UE�'��R��-/ImtR����'N}�ۃ��hf��ŝ�7|����r/mU����s�:�����Y���ǖ�V����=	�{x�C���;��LG9q��T������?���6�q�tt�(�W$�|F{�[�J �f���w�~�l�N�^�[��m c�Q�\:�P���6l1�} |)����F<aD��e ���fb� �w�I"V��I�Q�YG�� �98�k��J�im��)�ٔ?�3��'I��� ���OjT'k'����#��)(6f���� �����\˒e����
mDtc\��l��"�B6z�o"�[,�������?�Ў׸	�_J�y��;�l^ڼ!zb��+BlpjS��#ny�h�e�&�a�<���hJ�
��=�\W쥸M�oq4H��l�d=.:�eR�ZD�5�{?�38T�s��#Fϙ�X�Q*�uY����:�D�s7p��)%�k3��r�pT�|���;M�	��rgE�B���/���OQF������C8�ΨR���<���ObPJ�H���	xFJv.'\N�}tU�b(���NMP#�UM�f^��J2��8;*��S�}��Y�c����9��(�5e�/�Zc�3xR��~�TI��֩�n�Y0w�����K2熲�O���'������FW�����q_��_�lHJ�V��[�F�0qK�dk%$:N^#��w��B��Q��"IC�+ֽϟ*�R%�?�wU����)2�l���l�T,-a�y 'G��}SU4)7/h�OD?�HF���4� fo�>Ѽ���Qܕ>��i���uw,O��#��j=Q��ShI�[\(�I�����ߜ���S�\�R��GT�l�A�:�f�r*ݶ���ht�ah�Q�{�\V�2��`>UB?�8A��T�Ġ��O�I�X#�l�ü���L��A<Of��X��*�8�u�*���J��,���C/��5 A�f4�Xѧ���i��&�9�����:�r2i��I���4+}�Z��o�;����搞������Xɗ�/0t]��z%=8g���﵎��B�?&*+b�j,�T W�,��RUX���~R���Ҏ�wt� ��� ¾�|���z?��C�����򊽨�hn� �U�����	��sȺ�7}�\�og��*9P����o�q���o����#T������'H2��7�V���r2��;�����D�����N��*�.1��nEn9`l,�#�
�d�=������ωKI��/`�K3�G7���a@�R]�C��LI4$,���:�=��'7�ї�A�K�!��f�ޮ���
=����@*X�2:k�>re�W�U�Ϝ�E�$���)HԆ[$6~vS7_ɴ�6N�ش��,�����,�a���5y&c�el��,�
K��s�~:�B��E����`r���g��6����|S^�����X��{�L��W��,�y(���ˆ�w)
,GR)=P�C\���6�E�@�Ƞ�]�W(��e�?��3��Yh+Z���G �uC��qiW�pe>^w2�9!/6��Zl��Q?�4)��n�s���a+L�P�����]̌5b�䉇Xa^{�n��9~@��ɳ�B\p�@h���Q���_ᜁ��Bv 8V�-Q�'G`Đ~&{�sϣ�@��O�-�<��o�e׽ʂ��	K��5�-�,#s�6h?�HQ#p�̮�zhl1���(Y�^��S(NTu���ц�mx@͕#/5�/K�Uh9{t�<u9�G����PAnO�����Lv38C��ty�!��s(�f�<u"��\����H�οT���~���Z�D�%_��H䵘i��L:�=�?1�L��vp�����t� ˨���ASN�N[�j��u��3ܻU�y�+s����vY� V�\�!�M���Ehk���&~����e�Ɋ��\�l�>s��O�g�HG�����^VjX�����!��zK�!�W�Z�ChWG`o��KA<%I#Wۮ��1�+��E�ʞT���H/�ɚ�ĔG�Ʌ���geh�r0�fؗ�ɸ���T��L��w��M�R*) ���)\L�P��$�[�=�_�+���J�������a��󧧙N��A���.=�:\�"�W��s5��m�)�x�1-�(����=�d�h�r���cb�=�[��W�P�B�!)���DX�{�,�X����V4O��0�H��^�e乐�<�e���3�>!\� Ǡ#�(�������2�oX&-�礊�Hq�7��w6Y�����������A"c�J[-ԃ��F×lT\v"�!����ǶD��g�?�
~Ҭ��İ�����N��>s@:�� �`�D��hN����5��ayB!k�u���6��/r�zn�	&�`rk^�̶\l��qP��-�XV�9#�Ø�n�}�c
��̓��aI�Ge�m�5/g%]E���W�Z��TxۥeE\�p)��5]��RT��I!��R�$����8��HA�`;�+c�aˆ�:dT��#4=:vG�2E�b%@����in34���@BS�ήBtІ+�P��e	c>��c;ͦ�̉Ǣ��H:_�J�"�R�n���X��ߔ ֹ�d'��=?�ɯOZ"��(ȑ&P�m�-�v(늯�- �|Y���V��~����Z�����$E I%筸��V`cݕ+y6}N��Btw]Ұ��X��Ke@?/��DE�m�W�E��Ɵ���3��l8��s[@���ӗ�d���
�8��p�Z��0���mi�3�j7���4!w&��=ų7Õ��FXX��C�){ɢ�Lu}T��i�f]jz�}��c7\�sE��vjJ>V����Y�f�^�n
}+I�gz�!��F4�Uc+?�S���E�{���q���ya��M[�%�";|����?��^*�b�j����+��+��^f�e&7yK+�|N�/Y�� ���q<o��bmY�>�S͡vO�*����g�ߨdA�-
J�@�^y��8���L�y����5����>V���ԝe���ڴ�"����"[� �I�b�N3;h��|�4��$}N��<�զT��ﺶ�.����kD�p�u�Z�ٖ��U�U�?��U�*����^Ƞ��(��37�үR��V�Y���=��I�3��g���C�������H9K/mw-?6ʇ��c�����|ո�Ĝ���<*�F���?�j�`�6.D��!�?�X�0�򃡦
�����}��$e���jG��5����@�����t��-r����N�� 6��z���7�]1�[�˜a3�l��a��P������$s8QUՁ���\�Up�0����@�m|�I�����X6�0N`ݵj]�>
䎛1���%����dH�vc�H1�ʮ�<A�42�-�������6;�����\nΟ� ������+x&�p��\���B7{D!c!nކll��K�C�׏>f9xO��e#;����������_O2���#��<Y%(P�#v�tL���$�*�$�rĹ	U4��~���/�y/ʀd%�2���Rڕ������@���t��]�)��U�������y0'�ßC-�cM	�zbK�0���CP���
r���0�0�ST����ɓ�����$]��K|5�jE�wm�l�e�ң߂ �h����Ų%�;亓�#���&� �?��=�`{Y\�r����%l����Ф2���}z+ON-c^���\�ː����u!ըf�e_N�DU�y�݊*�)J@2"�]��a�nؽC��4uG�^]��������є�v��>w�'�z�]��33}6ӪJ�����m%DE���y�SN"h�f�|�$���dd��E
��(�WQ��A@�\�BwB�d0�օ9_0ã����=�o�]l_0%9UyӶx�Z�gdT H�Y�a�lf�p���#�������@H8�1�y�C����f Fﺡ���p����Ǉ���
��=m�����P��=eFEI�g�l[���'\���L"��xZ7L�u������vn���'����ʰ6��x ���;�r��gA>�� H�.� �a�C�"�)a�f9�2�O���Q��!������
6"�9sF��Ea���U.6�f���?z���V��9Se��R����-��_<����}S���P1Ϥ� ��q�J�[���Ժ��=}gq*�-�q܋1����w7��gk���<�������#�+���qF�n�gٿ�+A�1�j{6��h}d����D���܋����d�j�p�������ɢ������%,�`��/�iU���-�v>��Q�#��@��XP8���q��Ծ��}�x���<E��}�}�	�7�ne���ba�Os�0�,f/s�:�-��'��������Q%n͵���8f)����d����>�ook8�x�imrמ�4�D�R5�K䏱L����*q%��&�7V;�=���-x?,=>����m�]y��x�>G&w;=�����˼�	��l�rN
�6���� ���>�W^�P̶�'��U ��+�n��I�'�O�؛��٢8�+�o�RvR9�h�5�c
s�{���_��75�e�!���0��h��ۛ1��;����2��[����v�̻��g��Tkh�`D�.g�[��X	���h�u���c_<Պ�M���p�F͈��gV���9�	�����]Q������@���L���w�~�mr�����ơ�}���l��Z�sҽa�O��͵��/i���q��6l�A�{�[?@�o��@_B��>���\L3p#��/=E�p�G1�A�߸���&4i/�ނR,��{$�/z�$�E���'#2w�%�Ā�\l��ԣ�#�9�E���	�#a? ���s�;��Y�g�f��7v�Fbڗ Ktjɬ�8�eO`��o��0�JQ4�HB���3�Þmlbک��MCJ�:N��J3���p��/>Z��Rgr�ߓ�¬�w��̲�4q� �ԷI�.4r��rL�ǭW��>d�;j���1���F�ɄS&����L��s-	���6E� �d���`u�T߸&{9#݌����������ގ����TRh�
UE��+~���M`�_��?�O��ʑh�	��r�<��.��p)V{Kɛ�i2��f�r�(6F/�:P�ɼ�3�0��H`:�.������qlx.���*H5�z{��M*���M�3�CL���S�yI����b�%][�ʘ��FO(eHW��~)a�d�x�0�:��ྈ����Tv\�������(���?��i6�w�~]��������W�ƁXLލ���b�McӍ2W��[ܯי>�y����l���8*�@�����3$o�Y7�����J�I����>��!J�"���+��/^�d5k^h��cL�ai?Ņ�^��A�Q.8�B�:��M^U�H�}O�t�?K|_���`�~Ҟ�)x�W��޲�˚�<r�|9�(��<��O�?���>��b%Bc�%T+�yKa��7�L�gP��̆��n}��I�1��dM�u�Xٸ��,n�?���]?J�O(*J����g��x�Hj���9JqR��G�e^����JZ��jb��>�5�927o�mI-�̏�����ѓ:�K��X%�nߐ��?)&e	l�ӶTL��@O�;�Q������坒o�G9�Hv��'L.��36FHQ�󃱾�D��2='��m1 �����%�]-�m?@�١2}��'@�"��{�P
l�;v.���"�Q~�Q�&rF�"ȷ��ԡ�ݙ��"�ˢ�G�<��)vX�]NI�7����%Ȥ(�ڮ���n����Ң]�A���Y�-��m����U_�p�^��T%U\�Ԛ�qOHz�r7�!,Ac�5耯�J��������������i�AW�wAi>&}��3՟������d���~bq�FD^O���t]��l]*�+��*�r�p�G;Nm�ߖ��G`��?+)d�	��i�쇌�ޙލ�@,8jbO�e��F[l�5DɻNa���	x�!�����+�����y�h���e��7�O����������ɽ�G.~R��-#G�dQ{���`ڼ�9� ���"ÿ�hf- 2��"����u��kp�V��z��"�w»�� 1߳�)��A�!��?�;�:���؈�)X��h��
}�Grդd1&�S�����)��X��z�Ŋ�ΈN8d���n�.+!r����z<���8U'�S�Z�JO���#� �W�55���5sBNd�\\��\�_�tM?.�?r-!��V��(�Y��w?�ϛ _�l��B �Hg���d��Μ�{�c�h��\	C��'-��ĭ(�r; A�y�̿b�%����>u�_���4��Wöc%;%/M�g(c>�^��{�lC}b2ДL�2d�e���E�K/b�}I ��Sxe�s?â�J�bՑ��L���pQkbq����3���Bt��kD�HU�J�hg|����m�Fx	�,tE��g��V��c�����*"�w�h+b[�4�Q��HYw:I�Ӱ8eR����X��w���1b:���yRO���[�z�՝K�vH�5<�[�,��(~�C}�����J���R��a^�{a�s����䝺��0�S��'��o��ma�Q�]bB���,����.�Nr��v� ���/?s�7�����c�5ۜ;�N��ac�/\s	�z���+Z��:�.�)��8m!К��V�O_	�FvqT2���i8�6V��%�o}�����"��>�'m�}qp�����D�$[�Hs�=�H-l������)eZR��"��0�cs^�����Ty������pEq�Lt C�6�%�H4į,F��6�$&��spY�و�㈸MEBL��ѝF��F�u�#���w/L!+b�t���:_�\S�i�0�Y;�����&F��w[�dPr ��m{"Y�ۛ�~��)�Y ����&H�i�������375'���x����DH�����;0� $[Ȯo0����b=HF�:پ�N��~y�Xs���ʾ����;��?;���c�ޏ�����,�U9To,��{�F�4�yG-�h�a�'&�G���-�⾵�U�@�J�O�Zj�:@�p��6X׳��(/@h���N�1׎�6�c�mI~�����o���_,2�`��5᨝z�~��<Ds�'���r������@��F|�:�!����$�IĒ�1���t�������|�
���;�Av��IoO^��?����09�}Y�К����B�Z6��)q ���/U��$����297��D_��e�"G����tuJ�i��
?^�R����͸P�O�2��L B��o)R;Ed{~>)�w�i��?�[�Q���J�C��E
�r�k��ߤ�da�ka�{��0��<����Pc.�EI��)A�=
O*�$ �9��#f�DF�c��kZ��xL�����Z�q9aIm;���f�!�'KegѺ��pm�\�*%~?���]Q�K��ѫ�=��igt���2�����0aV�g[r@�rY� ��ڳ���q��F�a|�!ҟ�?3��Z*��Y/�;�	��YE�p�ega�ӿ���uvq8��(.h&�Z��qS��� �j�0b���Uq��L�>�c��l?�b�®���'�wJ�UL�" �n�J�F8�-�,()��90��Y��v���0@�P�~
7���󪷛�WƐ�c�(���1��%4��� ��V�����h��#4���B?�.��zS��^��0?l��N�5�?�8<��`@K�����}�*Fy�J�Ƥ3e�j����`��2��/~�����&(-��t���J���|���t�!IG��N�eO�����#�	�\�;-���r����z�s�ǻ���>�/6��3�edy�-럛�
�%����.���bg9�8��,��uhj��Y�5�g���Y<8�9���vfu��#��̄e�
�i�V�c��S��;L�'x�������d�w���]Y�鍚��|�6��3/گ$�k�1u�:9�ҍM�����}y"����Qo��b4ya�Է�S�:k���x�L�_A8�\҉������C��O"�b��Z�{���
�:Y�>��'���T⬿��tpp�����w�%Nw�?1����q�.x)&�!����Z>pʗ�x K��6��3�z����
�4�J@�8k��}3²|��W��U#�1��|�=^3���t��iώj=�<���b���w)�t(�e�Z,g>�	�ʢ�ӛ��a���C]h���e��a�p�~�߻�B�է��M� �q�Qa�$TY��m��M��܁���az0�i�1�@�T_�Y��%�	dR�q1�K�ݥ(���|g$/9>��L͸�$}����\jA8=�0� ���"r>(E��P,�ĕ9�Ft���@��v��抴��	���j�C#>�G�TT%h�#�ZB_Z�I;���	���g�-x��:�t��7����t����fw��AP}����CyL�6Ű�Tz��+H��d���hH�<K\�l|ۛ��M9��l�Q$�#�Z)��8�a�~���΂I7�5K�"�4j@�;���{�B,��q�q�	 �wZ'l����Ȩ}�W��ZB�z9z��f+��� x��u�lA�`ڶ=	$����R,���x���&�͛�Y��1�����8�_�|�=,�붖��7�.U�:�m�4�n�܎b�Q6hǾ�c�sҽH<��;1��<��p���Z��܇"����h��"48I ��l4l�j��v��z*�&
N.��%w���*��)�;ǵW�וԹ�tgDwXו��E�[p��
 �����H����4I�� ��g��֐�U_ ��	�>t�tzPv�pF����ܠ�����`�Ո��Q
���C>��q��U�5���$�[�QÒ�@�%[�3�l9�8Lt�H��U �󴔯S�=1KYg8D�Y�s�^�$�;}����[��oz��ڤ�M�+�[wF��/\����^Þ�f�J5/����Υ���\�����a/,�N�A1��0}2������s-��Q�n�;��o��Zr)^�2ѐ�_}�+~᪛^Fű��V�]q��$k�"�Oo�{�צgEC�6��R��va��i�ZB!��R�Ƈ*�H��\�����UPIzݬ�(�QW�o�0�������Ӯ���"�:�tT�S�R.�Y)|O�7��1�D1�322
p�Y �պ���o������-Ǡ!��@���wu��HV�ڽ��g���C�+ԂF�	�7�;��[��o���m�u5�b�b� Y�1���r����p�����y	����씪z�^��oh���k~�V�|��Ϗ�_@�0���~.$wO�ڤ���L��w�n����z�A_�?�-�)��֑
l��;��Ju� �;��
�h){e�����9�u�V����c��dv��c5�uF�tD�L�c{MX�����������5y�m[�s�c���l�(���
�f�L����<k���sD^�iᡫn�u�r���˖�ω7	�1���ȡw2��ns�����xŐE����x&��;"Sԃ��f�@�t�vMV-+����+�Ʉ��v��y�����;sӾ�Vp�RM泯E���&�鼥c�E��Ύ��>n���Qj#qg"z��7�R�1��O/`Z��E�����M��J4VA"(a=Eb6�U�P���7j��PR�����7xd��w���v(�yVh��F���1�ߐd�B������	���>�ɽ�D�fq�o�fm��*����_�4� �t�5��U�,�j�	�E�1�U�h�_0	��|��d�,[�=��O�o��j&d2h�4�����^/,���c͉���ʂb`d����$Ki���ڽ!���^��6��6�E�����49������L�qD ՙ���]8��h��$,��!:���8��R��������+�vp�� GE�j�cG�Oƫ��Cv�����'�Qp7��g&�J@�Q��!E��)�\ʴ�uh�Ԙh��qJ�"�hS����\N~Rg1���}��E��V��9^�3w��7�*�=/)��v$]�4�mÓn�*B��C:~�P�[ҠR,o�(6h늺_��=ojP�՝�9OS�A�pk�_��n�D�Ց'���E[C���2}��@�A�KE@2���~��M0eGcⅠz7L��&I9Ӽ���c7Y��1E_d��V`��P?�&�6�E���֊�Y�����;�~���������q]Q#��뼑�+!���hki�:A��=����<`�5���-�G�"B{���o�}2���E����?*�0����*���P�t��mG�2�2�M�t�YGc��İ)���?�>��!5)W%�u$y�ps�����s2���pU��imA���94��S��p�B�B�/��dCjV�6�#��%X�78&��UBvWo��H=F���,A܎�Fo�yw�X��K���[c��68!�p��@:>fk����a��LC����J�&�ڑ~��̡�V�\ ��5��% 9U�!@�@[`,��a^�k"�m�A��{epJd�br��S?�4��4��/�ǯ��Yx�e8�Sy��!��A/<�H�?KD湍�~C�<�pKxSN-A.�46�@�ʚ0" GZo!�C���ЬF	q�pb�ٹT�c�o!�ˎ�hq|pcc�oR�A���O(����|�w���!���!W����ʃ&�G:r����,��5����?�20gM��_e����6k/O���|G'��������~#�a4����
��	�t+��A�����T|F�3D����\�@�O͢P�J��6��uBJ��>4b2�&B������;#�E�5�F�����aYS��aӂ��G����\�!�y�$�'W�gRa��+]�&�w6�t�'3\8B�{(�u��X�����y�ƀ��k���j�|�P�#��y��{�$)�<ݫ��dG*7�+�d,�r��t �E �kqI@�I.�[뵦N?=��I����:�r�q�C�ɬ?��^iK�f�L�R�R(Ƥ<�_�f�|b��K&(��E��-0c{�Š�B���+6V��+M���O\�b���+�c�!�]+U PIgz�❝�C?~�T�G�)Q<W��9�Ԉ��A����?z6]iWֹ���G>S�y{��׶���r4��b��f} �t�k#(�gpG���r ��Y�j��@�F�SǙ��7�x�B�����{Z��uM-qJ�ފ�b0������<�m �5�Lx�U|{`J y2�����Q�(ȇ�J��y�Dw���B-��xr�ة��v/���x��p�A@�j1����iV�����|Tc��g��^�Ȳ�Vc�q��X���0�c>}W����&ݢ����\�q�"7f\��,�cG-B-�􄱛��H��1��eΑ��Z���G"0����A��p�S�c��}���35EK�ga�Sod���nek�Zl<�,_q�PG��;`���XX1��hg��cw-���}%NXZ�Qb����I4���1�BJ�
�,��U1Zq���n�3#*�>��V��Ѽ␵��ȲΡ�$��w�7�-�5���C1L ��A\9���:Ҍ8�w��i�M7΃��K��{�<�%jL���h���.r���P�BC�!Ž��t��l ��Qp�v�:c��%$���3��x1���.���cȏSq���$�0��	��\��ޥ��E#�dIT�6���*���N���z�����.�K�mY�yk��9M�Qi�  �Ȳ@��k�V��㏀ǁrj�3�d�`���� �ҿZ���?�*�١i!�ͽ8 �RO�M	#�PL�_�n	\�䁰L5Et$>k�ޕ�q}��kVS�>@�����m��f�(�7���]����9��N�xT|�)q9�t������n�=�9=�L��I����N�leI�Uf�'>�B��F����O0S��������tB͙�
�m��r����W�'ny�h{ڮ]��|��*X݀#`��e\=��W��k^�o�G�ߑ��(Rw��L�<s������/K;�$?�<{�a}�d�x�:���}��shſ�ݱ�1���8����6u䀝��h�m��LW+`��$�FC���A	��WC�����nLV��S_���C��I�O��ǭ��\	#�9c2��T#����8�P����u:`p=3>����nt4���5�6D<H�҇-�Q��0���G���N˺���>�&��!e��C��N���Es��C��Z���
�i5p�Bnбʒ��"MݧUq�e��C�2#x���q_�+?�O���mawc�XT4X�$��^Y��r��[�z�[�,�h�����-�ι����&��L�}�?�R�0i�<uump"�R�b��Y��Q8�
�L8DՈc�S���D�\-���Y�)��3��1��9���~C��[��Z�BL��?<ce�=5�\4�TJ�Jj�*0<����(�s�2�?Ř�J��ut77]��Ӿݐ,:���6�"$� o"���Jގ��c�4*�h����H��H�7� ��I���"���^(�4��:y���q,��~Hk� �`�����!0��\WHΎ�*�K�@8�[P���v+�_��vD_	u�F�Zk�6Ѳ �<$�dۢ��3��y{�Q�
l����۴M����1d�*�!Q��_���{.x�5��h�D����j
�x��g�b �$s^�(Tn\
��l�,��8� �ͼ��CF�nrr{[��S�/��V}͆�p��<��~��ڎb�-3�óX#=�|Ƶ�wR	���Ќq�5��H_>��aѤDr*�A-M�,�v3��C,��eT�0z��N����@`me�M(�YE@V[Q�-�V�P	,��g�p1��1G����ە�a��9�2�X� ,ֽ�KoRip�6�Չ������A�/ө���Ǚv4�=&�� :#akf�g���)T���GJn]B��S�'_����3��]0�fM��՛��I��ŏ����2Z�J�5��_�O�m�֌M�� w�F�e�wOT�~�/}�����UM���8��v��j��|������������i�f��c����3'T��ᒲ�
��'S*Ii�;�	��О����������&�d���%����C -�����z�Z
T��ȁ������N�┶%��/A�Xj�4��=ՠ%�� .L����_iD o�$o8��{�'@��@֌����7��5O�KQ� !�
+lҌ��I�KH(�k����7��{I��׸�D�t��x���u��f��*&&�k;y%�۲ �E��2M���"Y@� ��IvK�iy�`,�c��G��ޓrR};:}J��h�P�ќ���M�*l�fQ �=�Ÿ�- 4�M7y%š�ul����S�Sɠ��m_[���D;�>��+(�B��
jr���wU�!"p����Si�������K
CW�u����
P4Gz;Q'`1�j Cq�iR�^�1DP�\�8�9�еv�0�|J��_���׮ܦ�WO5�C�춘����QFi���7Y
��!����]#�!+�	:�m~�}k���(��?���qu�>SK�&�\6���Z���OOa�X����{F��5�B��1���t+a���7�O��v��3�BM�X�D�v^�"������%)�g��`�<�4v�g�	��%M#�P1�^ 4�Q&��W�V��n�������=UK�GK969e��ӥ֞b&oY��V�!�����_ZXٹoIF��Ĝ�\��8E�(Td�IЇ���Y����O��ip�c^f � A�nP�6l;��B
$��Ut`z��l�̦�n#}:�BI��'>%�������o��L|��a�7���L谊GL��i���oZ�z�W����(j��;v�6K�Mi״s/N=AZ�/�&��3�̋-�!��6��xʹ�3�-n��5=�?7U"�5�f�5>��!@�CQ�]xy�����ܐ�D/)�eW9����}���o����xD����ww`��bFU �|~Y���-��ofC.�_R�M�2m.�|(E��F���s�0Y�*�m��]]�����)��Gq@2�g������b�Tl��B�m"��X�Ę�C�&��q�AG1�"ݝ�]e�U���,a�1����-����-��/ Hw�9���Zق�@���>�H�"<�"�����\.X�O�z��\�N9�S�D�~c!`�T&��?��tzpίAW�>�?�0'�<�:�}���pu���|��c&���Ȕ��f����[lbT�$Y�:U!�=u/'9�����RȿAN�W1J�E+:qB�xCߩr��C�[`rt^�s�����+�e��̔)+����Ko^�uy�^���F$���M��p|��>$}�ɤ�۩�D�o���v�A�� .��������|}y���X��Gh�%���C����~�\s���-����������ui&|�V��5	e�+�-�j�`�n�QS6�e���Z�FAK6ipS3��1!����a�;(�ᇽ�،N�)�%ws>����o]9�f.p�O�����Ùs���i���mXLWV����MM��8o ����O�p�x�i\�F��_�7���n��L�7ѽ!ꥄ�;
Qa���/��r�^�I� ����W��X9�Ţ�o	�.A`}D��Đ�ֈn)�R�L�ܷ M�(?�;�~�ˀ���bZ@��w��3�b�����(jx���cdG��NX���gzW��G%K�����,Og�np�ĵd+k�=�������w���+��_�1�y�'�EG��IZ&���us�y���!Ww`���WV��A_[d@���9o.�R�s:� B}�(J�U�0�� ������0Ɍ�1��{:A��;�t�=�2d>p��ۙI��G�A�U�����RD/Ǧ3��,:�;Ii_���za��)��:A�T�en@yÞ\��+�a	h|u"�u� kQ�9�~0$$	t��iL�Å.�G�m��C|�ep]��EYr�2��+��L_:Q�+.P�޶}��UI�3U�xp�r�9��bQ�z�:`Rؖ����o�ֶv�G� ����	�?l�+a�,��Zx�-����&���GZ�H�牀��>�W�)K�Y|M��Y�6������Z��݂�|������F1��|'�.9+x�}w�E��E�1A6U�U+Ѳ���`Y��F��5H����ug��#i?v��mɉd���~�Z]�S���O���JD��k8ga5�
s81�^+W�.
@��0��!���π1���M�Z5ӏ�)��A��VI4�LW���RS�U����H穟a��aTY*.���^uB�����{0S��G������v��4 ss��+{m2��K�:p0�I:�wʶ2�h'��*!�D���1(�T�C��`j��eW亱T)�h��Wif,�NAh^�j<z�:%Ѭ�������g�SY�[IU3�@��؛��&'P<;��rڮ�[=�%�i���C��ސ+�ǅ��ΐ7��Ɖ�8g�Z;u1�h�`"�W��_�M����������%��@W��d󕚴S,^�}I3��y�D<�j��6�/l�_�ʑ�]l�v3������kMh���0M��<X�+"�F����Gr�yӹ.,i��f"������ fn�b�fw>���%A!1_G�k]� d�DZg���N�?ח��%�w��ӥ;w'�(p}Zg�������NZ�@!�9eVE�pXB0a?;�&��q��<�t+�:�P��hʰ�v��=�NQe3� "���o2� ,-�P�Pt��v��A�$%r2��m��u]΄�ݳg��~����A6;waheN{tw�k-V넛J����j2|o�c��[��b����0���B���<��.�M�q<�/�l~�-Mn GK^hӸ�!��������c����9�k�y���cL�
�luH�+��tj�Sׅ'l>2��e�������+~�7b���d��_�T��_�n=�m7������m0���U�2l>�HE[�g�A��x����o�Ə�q>��0�)G��B�7���E��O���N�Ͷ�Wu��dIz�x���oR��@㔷���\%V$�^�O�"2V�ú0���Q̎���][6�?�L�F"bZ:��	�g�Y�3y��)JԨ��9�1�+ 
���J8�g�cM$6ϸʷ�]S�^��H�{��{��5DQ7t�A�^'�@`n�|:�7�lu��������n�t�����y�58��\�[��`�Q�F/S�z���7猳��w#�;D=R e�	l"9��z�����I�uH)��ôt��b��
� )�W1&��p���4��Q��q�';g�#����BNB���ր:� ^�Rܤw0�.�A/iy}��Q`C�}���8�J�_ގ���U�8Z�)L!�=��T�t�!ό�T6�P��z|�x*[>$�q��>�$���膎Ų	I}���M�8��Ak����`#"�]1NI˻P�#��U�M}43bR�KK�bT��])�?s�7�b�ۓ5���a �dA���N�ڑ/PA�3������B<μ��m��:�֤4��PE�̍T����abw�^��靖����T༬ym�$�e@���y �)�&j8(�w�A��;�j?�̄��-�-M��' �a�J�1^$�Cqq�i^��Ĵ�`@�?nl�1:O���) ۂ~���=�/�Pp�8چ�?eM�߭�Β*��܃�5�WX˷�8yAÕ�4�΍tqՁ���K���,ƥ4ԕ���,�1 {�(_�jt�N�j��Z�cK�ru�ۭ�zRMk����Ih�Rd*� � ���n@&տ�ۑ\G[�l 3�D+i��% W4^�����|CHww�AyȰ.��|W��)�rw��( (cr'ءpvܠ<[b��<�	��Ek�T����~�o=� @�~~�i��g8e�T㲄�+*#J:d`��e��DN	�3���Yޟy��(��nf-l��+��*7x�$��[�NvRµ%j�~����1�+5cv�7����o���B�=DfڦM��j�j�yjղ�#��u���J�[=�ի��Z&_����l����=M��rZ����o�Q�%�˨����H�+�Z:�zfy�1�¨���a�[��:���"�%��2��/Nm�-��wQ0#����J�a�8�"��f�ϬH*�D���ȵ�eȄ�ۮ^&:4�ߔw�Ƹy�/��R��l����O_x���'-5ׁ��%Y��̛D�F>.X��ׄ�|Q�/��� ��C��C�l �ض�&Bp'�����	�烗�/A���:�J��	�{�K�?�����tR�7A�(��yR�v=���UFY`�MoZ�V�̠�!X�� ;����m�� �/-+u~�؋_�)9�nT���3�z8Q^��Z�8N/�?��U�.穔u˴M��H�*��	����!�Z}^+j���?_]��3k��'A�y�ռݐ�xw�Y��\��n4#��7]�Sîe�Y�i��8\ ���7�yeުw��ә�� �CT�їVt���z��'Y��}����p0l�(�����C��L{���U�X|ZG�0�2_�5�"�>޴@��y1��C��j��o_iF�x�yx2���H��]�2�!�$#L^G�t��ܡ�b�P����[����he{=�@E0�;w� ���Pj����+���~��k��T�V��U�mz�׷�x"�j���V�@�^�7����h�����=8�a,*�+��/�^�Z(q~k��;�'MT�Ws�"����nPdgC3��OR'����U���訟Ȏ$�j�?$���$ٺ?�g y:��T3����(�w�)�V�h�n}?���.��%��ܞi@�o%��x�Y��_N-��{cv-:��[@:+W���ZY�����Y!����K�����&8*c]I����>H,2�o��^���o���iz4��)xTs+��_���J��%쫒w坨J<p��P;H��w�����/��Q��c#XUUzd�5��wH��]�x:�<�=n��9�t5�D=4�d�L.W��&)�|d�9ԣ�l�&�"�gr����D쎙w�c����C��^�$�'E,��D͢�8͖��b%!�:d:��oQ�UU"����3��\t��1�9�~�B�� ��,��iv0'1�cH��_��_LZd������I�eܴ%	��˯=��O�! ���6�/� �~��:�G1Z[����띱-�4%��0܀k�l�z�~�����K��q%e��ж+��ߘېP���E�����ۤ-���5��*����T/��P�1�;F�X�*��~�g���2����GӞ���_�c�¬V73Ɩ���
2h�C�o��0
7>�R��r�$0����i�1��I??�L���U����p�̕2v-k��g6��?VZѷO���rXH��oo˽�TG�.�`���v=;�'���)���CC�f���5f,��))\���<[{�'?Oc�v2Ҁ�}��ۆ,�f�@_�P��sa����>$�쌸���:�P��s�G������M�xئj6
2���Z����
)G��;��e̰�����ϠE��F�%Yt�`9�|1�ղ���2�;TK�r�y#��_���"��0�*٠C���"��	�#ΏV��Ď4a1eIh��Jt�������(��tGn�;�[C2*uXr�7[?��R� 7������ϼ ��Asz�F�%�hLq<#'���Z�ҩ���=�y8s��{xǙq
���u�A�Q0�{�
O)u@�՝���G�bu�i���E%F�'��m˯����K�&^
��P��g*�i525+h|�R&��طD_��0�`�,�i�Y]�{0\�����8p=�ZR��e���yK��E4	�7�?f9�t5@��ۍ�]����e�z^�w�b':@�=���d�+�ol�t�)�)�o����o��֭�S�� .�;��\�+���&cÙ���� �$�~3�櫜�a��g�L����F7�7E�&��ծ��� >���m$*D�CꞬ����yNg��]�?��ROk<�ӌ���k�9�Z�ʶ��8���k��+o��Fa��������OS5�n��/�s�N�����d�)M1�Mwu`حg��V�If�F����e/�MG��1bhmK��$�����=�&}��uJ!���u�B�6�����r�q��I�V�2�ܴ���/��1�g�����*���*��8�m�����:N:�z�O�O$<���k����>a��8�s�������F�D�S��\�Q?��O�1r�zf`U�@JM��{;O��M�s��Ю۸�5	|g�7��6zo�*��Qi��h��ۉ�ö�2�� ����♵1���@壶�אJL�1cV���>�+���L�Z�f�/�_jX\8#q7�^i@�̫r��D��a�<cH2�*b_�]o�}�����
�5ocj���P�)��y#z5nl������K��bbHf=��7zHL\��Ň�XV�&Ң�I�TN+�x_Y}����}W$F�u�Q�"�cx�]�1>�~�3�,~�� �����cY�h p�j�$�S��=lL�+V6-*��b�u! M��c�<�V��{��P(��o�+�2���"�j8|��jZ��y����x����b`}��f\b���w���Y��aW1���m������LZ��_��8n�-�턵�l���]��;�qۇ�y�K�\q	�X,�m�@�8�\��<��߀��/o�(���O^"�M���R���_�R��{�D�t�Z����!�2Q7� ��Μ�-l�a�?���\��<����߀��Ԋ�߰��΢t3�EAL���>L��r���M|&@	�8���������x��8�	�>R���&�.moG��O��:�P��>�c�+�ߏUV�|�6|��2���JDCV����4�,^���ɣ�߇u�m�e��i�B�F�e�şmH�1K��o4��dRI}z,Ų~.���'Y��Y�de��wx�]_�A�`鳙�Gɝ�#�����q��7h��]�W�2��ًuuG����B-Xx�����ײݛ���	�����b�������Sr�2Z)����گ;M�}�v��k�|t��oL s�H��Y�:��N%d��X,���.���F�6�;vGC��̉6�\
!.�7�����qs�����@��Ol��Zi I|��}��cSo�v'޳e@ɇK�Oلz<�Fp0��� �m2�B]�*�%l�(#t�3a L`��v�G҆����x�ys��6��AX�<�_Ry(���7o�0�sG7Z�_��Sc0�h��oC���#%�h���Nf"��Y�!3�t�`���k�z^cr���F Q 3}�!��Ə���z?��`�IaK*�Ma7��>���K��dSP�5N��lW8�|��{J>�U�lT�Qܚ���Y�(�8�>���i��X0�R|E�&%�zXҗd���4\��em��;w#&̖A�"���jR!x���FA9���zܠ�-�jA��6���[��B��=m��B����o]J#��JFi�7#eE%r�4s̋v[���.���m��o��O��(p8����dj�
sm�=C���Ɏ��Ȳ��F�j�v����r~�=db�x3c�t���/%
�����c1�Y��Ν�7x����u�mVy�=�U���/�IDu���0�.�^#��sR[��.4��►���b$m�)MR�dy��J�ݏj~��δP<��ظlq��^Ec�����ת3��dL�'�2 x�OZi���t�4��'�K���S_5(����K+�\�2xf�&Ɛ$�")�Fs����z��T��?��w�*�?9`�0�f֋�`�8�x��@B�u(��]ڮg�\���k�R�RR-]%$2�bV�)k "�ұm̗��qOX�a��!Ɛ�ů$�(�+2ЪRq=1�)���Zx��dv��#'}V�cN��[�߷�Z��.��SY9�1��"�t6stme^קXj\��#�[
�� ���<W	[#X�v���?ݿK�a���ߐ1u�Ґ�_�!�o�yޅ��%�CE�
�L�p��ϟ�k�"�/� h����o�<dH=����*�N��ej�=�=)�:u�`��ec���^�p [�da�$�.��:y�uD:xx�yQ����X��O�\Hxn����j�`|D��G�,���3��R��
�^�r�K���	 (i��)WW2�����X�I�ݧ�߽Il��ߌ���v<�!�x2�7��'"�g�JKR��'��P�D`�a�q���]����L=X�M�P����^�k�<�F>���`m�����d�x� B<4� �a�XFy�[:#�����X7����>�����7$��lj�p��"��m�������O3��#�����a��QY�;�����֔�w���i=f݃q,�P��l#��3�q-���w!��S�t���7	[���
��[� �ʳ#���;�&�v�w�#�@����X=	{+����VyQ>��E�k[x�G����Z<�j�'��n��pa��{�uKf���F;Z�ꕻi���u�����H�ӟ�ӓ�֟�i��K���r�l�yȒ}�ds��t���3���a<�~�����E��b�y���P����L�����r�s �)F��PX���Ƅ�*L�9pS�h�vD����!W�.s�7��I�H����'�U�L�y6����N�Zi���;�aB�n�h�y$�:[)T[|�F�s:��!�]�S�|�H��8x*�z8�F�6k\or)�!��ߒ>Qo?�������ɂ���"N,Ž����Xʚl�Յ�.m�Sz�7��YO(8��Y�B'��d�݀�����-!r �K�DO�j\[�o�����;�*K@Yg�� 8������-��ލ�֛�^	1�Д:��# ����°�����~ �{�!����N] p����rqȭ��?���Ch�Ay�@����пY�<wX�õ��Ϣ���M$�?�_`�	Q��+��y�:��GV�B�<�y����Sr��Ե7Z�H7�l����{Wi�W�����B;�<�9�C
^��.X����\\2��VڐЄ�k"d^�����|=�D�d��;b�!�LK�V��w�|).v
�\��m�#�p��h���:�Zi����o2��D�%1���\�j$��>D�gB�?ko�|�@�f�W]��>%�bx����5�Q����xM+����2�a:T1��	�5���M6s�� ��(�S )�~�w��"N����;��;���kd���nޥG1i��1qc�`[����B~���jEzu��W����b���o.�����̜t��E�x���I�������U��b���S]�����k6���M��������}��
��sh�������e�
Q��d��d>�������&��C��@�����t".��p�!PNqT����=t
���.�saShP�o�dS6�3ݢ2J`x���k��/�_Y�n<b���k�4�^�ŨR��F��w�p�^����ư.�7@�d��$�����e:P��5Uu����m�o_-Pz�d��84ڡ�o+�LRnL��m� \��mN�ǟ����e�ƺ�LM���ҒN�e2�E�a ɩ�͝�N�7��cX��������3<��Eb�:Va��v�`�*�9���� 4��QɃ�ʔ5P]�����iS��L�m�kg��J���	6F4��!�[�%d�_�_[�3$^Ϣk�f*����Sx,c9Eq���ܬ7,��|X�;Bk�&�6�Mt�˲>����{���g����k Կi��7�Y���J�謢=I�O����+zU�Yd7p��m �O:\��3�?c�- Jdv��QCq��&.�.E�=QR��^ƃw�8D�Y#Xs�������3Ǵ׵�:�^{�c�=�������CG↦(!�DK{�¯�Me�=L���ػ�}q���#�N��W|I7"��3g��� �C"9��!�ԱC}��ICh�7Jq�$���[�m�!k����YD�H����ǁ��Z"nQ�k��������H��fp�3����B,ݐ�߼�ΐ�[�f�����We�Z(_ˇ ���q6�����*�h�xį�B��9t����	"�c�08�}cY��\�`����#K��S&@�~�B֌�`��������v͞Y����
�l)mк\�������s�0�Άs����2�Bכj����!Ba�)�b��8� ]Sӵ�{���O��S�fj7@&F�M;�14b��&��x�*PAYf%�w�>6B�xͿ�����1M¡`�5-�=��}eT#n�Ԛ]L�Ff@E�ⶇ��C�U���=9�̹����j�������*�xMf#'fi���S
齂"<�wA���f)_����K��X
����{���C���.�n$c���UX��q��
��8�x	 C��K�����!9��mvÓCz��#WD�� g�:��n�'D��?<��#$�ٲ]��&��sV�E�Y`�i���� Y�-�Z��:�Ȼ5!��)�էt�CY\yc�q�+��\O��Hh���g�j��c=5��Kx(P�E��{����J���.;����A����~	��d
���Md�Ϝyq�;Au�x<��lE�����Q���q������/pf�t1�Ȏ�+Y~r���_[y>+�7���,�tU�9O��yQ���7_:�M��gRk�*��F�;�\�O+�n�^S��򽌳��_@�݃q0}E�8|#}�I�vеc�Q�C�A`�݋B�ǋnVަ��%�-ʫf�H�+��`���	_��p��v2��3T[$�(y��B0[��
E����1�w�����CĆ"�гW$�=��'H>���Yee�p-({v ���´�v蜫+�}�ݞ�Q^s��0�T��d�:�{��3�M^�[p�6>�(�ʜ8�y�b�/1���8reƆ�̃pc�ͅ޹Mb2����
�X�K���S�QW���+-��q��X��\�JF-H=ƺ��.��;��je94�Y��/�}�������n����ߜ����B��^q�y��s��Yi�PF� aU0��H7���/"�Ø���7ثԓ����WB
z&_��
�W���]̈�kf�5��za���ШD_�Q%{mx�Q�Y�`o�|}�����/��j�]�8�۩tf�J�©��G�/���<g�]g˅TUM���'Rr_���~7�+:C��r���z���a�z& L�B95�1N��0�@�MM�<0�k0ϟ5[6�rLq�3Q�T
�����'_r�����y'Zj�aw,s�$Q��t]�E��.�kZ.�[�;�D:�^jg�E=�9��"�.�U%�G͟^�b��P-�Ⱥ�Tc��S��h�f�0#���J������%���>w+,:�����Q��I�pN�?�h�9�l:��r&���>��]x�A�Țc$S����S��L}��`ٓ�NA�T=��lo�XnYo�Ui��(n��{ԕN4^Ǌ����4��N�Y�/���a nl�E	�3��7o,/��K$��E�O�P�Ze�۞�)@NWtMt��~�n<`D�[�BV�{D�Mv D�Z�|��l�8�f0��N�����'� �w@B,�"if���S�чL�F!j�շM���&(��ĩe�r­�\E��5�
�"���/�ɇԴ��^�O9�4�7�r�{w�"X���J�L��]"��)]钲�KJ�� W������;%�Kķ^|�4�h!��]kղ�\�.ȿc� �qi���;圕{��co�i�v)�p5J �\�	S��N_X�i��ڼ�ܭ:5���㌷��童"&�CK��L&G��V�f���ZU�;1f0���B��ڑ�>J��`���o{	���e�o���-,�9��$�)Y�c���9kjA�?F��;E��x�_� �x.�N����l-��H�ؠ\���w�#��C�J@��Y]l����g�$�=��� �-�P�b;ED�9\�<!�E�ڥyη�`J�O����Lcu+-�J��Z[@��GcWiW�WA�����A�X�Σ��$����hƮ��h���q��i�\�f�(f]���>~��eKÍh�Ke��i<���wmlB�;�}��N3�,���i����A$�{�������em.�1��:��]�2M�(o�"����P&�"��Y�{VH�N���)D|(��M��>}*����fx�@;�Eѱ��j 0S��wmG��F"��:-�6<1��x������ZI$�A����&!e4��Ws�R�e�l�V����Y�T��ZWI��#wL�g�U�{�a1���������w��s��H���Қ/���3�qwz��h#*|�ɮ���W&owu��Ie�C$�B?�<�+��~������MUV'�C􇜂�"�rW��-����AhKfF^cV�
�S�W��/G�V"��q�w}�y��6��&���s�^�HzG[&'E6h-�(ZO��N��:KT� ʂ���ҙ���n�3L� \����:��R��3'�����/Ԋ�.�(���m�8��j ��<�݊��Ic�  ��2��a��a}7�m��+h��VA���+�CYƊ~��%��lśjd�X9��B��(xƅ?|�ذ�gy녷�գ�������z�#�u��\9Ѫt�~e����P�_,�S����u��@���E���-*��D��ζ��{�L8g��Xfn7lk�%-Z(j��bxYy�b�~߇�um�SEϠä*#�HgN���T��45i�~� ��g�:7���'#��ơ^���������r�C���.[g�le-v0Mk!k��26ՍHt�j��Д�?��>g����LL���Z�߫��{g�E������Ɂ�%g�SRM��s����)��	����/�,�����Ư�8'^�5�w0����!�d����;(���0Bd�Vi:|��xtn=���1�P�P�d��f	L|������LELaH�:{�ȦtU9�-�%06��nQu���9���X��xemB=���5k7�x*�;J\�Q��x�`�Ľ��5�-ſ�=ٺ�ד{�?D�b<�~�?�B� ��̈́h�>Sdj�D_���Ek�� ���j��;�a�'�Aہ����<J6����Z$7 >�ގ��q7�����+�} @�}�,����զ_f�?��:?�B���KAPZ|o�ؒx��>H�u��צIL��������|#�!�Hf�{��������Bo�����;����̹|f�ȼ�ׂ"���9]���gK�><=G�<ޅ�'a�߇+Y�)�ג�ewhP���~m9{�r�{?c|8���Ӵ�h>Ql4�G����|�)[�X��@O�nZ�~le�#�O����A����K�����$�z��Qs�>5�MW����8�%as�Þ��3"g9�nJ.��皒d�B֊� �*\_Ze���@d��}��ya���}՗$4C�	3����ӈ{�J-����Sǯl:CZ�)�s'�uq��3�����?R��-:^����N�ҝ��{^0���i:@Mؑ�ܵI���9IO�Q?��@��v��zu����-����r[y*b�3�8B�ܛ(a���H��j"YܖL�3��'�U~1)&�M[�J~*��ӈ�-��5���>e�ww�i���"�sQT�ٻs�W�x*#ߵ�~.�P��\�6����~��-��e�R�]OJ�V����IL�fe�.�:Ga⶚޴b
���l1.���oĹ-rpG�K����%��Y�~{l���u�&��g�c�0_�7־g�'~p3d�(Z�e���"��$� Ƭ�`c��3��W|�1�T���IDU>y����ʓlɠn|+�^�ƞ��qq'5�o]�k�vW�شaw��d�qs�i� ��0�����g�!��<���ws�|�>�%��+Z�ӆ;S��ғA��������U_�h�87-X�B��jE�z�ӗ��zFqג�2&5.�u$2AM;c�ͺ俤1�"	��J�VI�#�z~��l���G�T{�ªB)o��iZ�(���l��B"L��������ܹ�L�khJ�~XI��H�6�F���s 8�UҙU^�EIN�Y�:�|���S��U2`��6��(�=��B�A���u�1N�^�����β��<P赂�so`s�,HN|Ӹ��k��$sվj����WVbҗi���Cz���6:�-�`K%r�e{�*껮K��۹�V�?vR�8>�rf� �<��5
��	��P�,aM��B2� ��uV�+$�!�*\��*r�*�;�✫� �ī�t'F2�g�
QG4�H������������e`2"^�߄8��m��xTVU��kb\ݿ٘����0�B`�ȯ]M'y��Uy{�-����H�9�V.4��)�z��FC��³�ը�s�M��Uّ�ϋ��k�0�`rI�Wf�����;�oo`����E��k�[�;�{ i���Uq��)§!��Z��K`�:3�2��|���7�h��@5����K��%�c���@�����o��gj!s�TL�{���>�-x�!�Gw�bO��Qc�o"e7_z�ы?
��33�8"i��H�1�ĄU՘,��,2+�ҚU��*�K�`T����r���)6꩜;���>C���h�ӟ7��^?t�"�A�V)��o1�H����3�-ς�]z�r�e|�e���Z�C�J��3riX�R�u*X��Tݩ�,�S�P��>�Tx��ؚt�P5��c����3��21(̡���2��^�QX'j�b��w�  ��w­��U��ˢ7-۟yEW$O�DE��X�ݠ	�D�<*� l�+�n�.��X��3ӯ!_�y&Դ�9ѕ��d7+Zyc���#Y���?��W�|��\����j� b�IJ�C!����n�J ��S�:m',e�&Xc��B�oe�3M����I����ARb��`aF�v��h��}rQb'�*�Z��Ҙ��_ r9E+�ߔ]a��m����9�L��1�?;��Z����\H~I���nxmP���2��J �$	@��9�����R��=z*���1���l��� u��r��ѳê�Gx�y�8H�;�	�b��; �����Y�=�Gȷ4�h�z��C�l�m�����8 �}"WN@�:k��3�|�k?舏�y ,-�-��G�a���Od��e��E���m $W)q�q6*�Yx��4#�2"m�2j��y^� �;��F\�\>v������C�x�wJ?ʂ�����yE
�p���w\D�7��*�M�^3@�o�i�J�W�y�&���VFh�78s|-�;N�� U�SCン�=��v7�!�U�v�Pa���&@D��љ�
W:)�>�ͬ89>�t�?���{S`���v@���܉7�� [��ӥ�����X�WU�DF�+��el�F_>f��N �z��\��������H���F�il���j�c�!���Ô3ڕb����1���W'Oz�*hc�N����Y��	?|�ҍ�]� j�z�����YI��e��62� B�����5���`�5��N��P�rg
c�T��fe��v2�[OП��_\��K)*�%��C��"�Z+�2BP���O�Z�(rŞ��q��I#m���܃���3��+R�����ҨmK����o��:�뎴6������Ojk��%ܶݱ��&��Q0ہl5�)rW�]B�UZ�IYh��\�U��h�z=`�'b��Ц�6�I0n��_���k<Q�����E��7i�CK#���Q��q/na|�Axo߲�p2�Vw<?ǼE<W��i[=�+���2���v���.<t�����zO��Xd��C�e�Ge���˰�!���r�~�E�Ϝ�t�('9@aL&�<�Y��1]��pRњq����<��wn���U�,�r��y��Y8	E�FY%JhgN;��v�y�ɨ�17�GJ�����P��?5tlw,��s|��?��W|�NGv{`\�m'ѲS����|��j�R`J�D���Z��p�-�]@��M 0+P�,�O�Z��a��0�yɺ�Pq�F�mn�+����%%arU�u��6�r\6������!�do�4{��=���r�e�a�6_R�9���cR7��p��x������< ��n�Ћ�ncg�wR;���@��Wεi����.u�����m�BlY;�-F~�'��u�[�3L��y�n�=^`�
��xBP�������6CM^���������b��*eį-&���v���|��)���H%����1�r����F'�C~� ��]�-�-�1Gى��}��&�=Qj<:O<�S�T�Cj���Pn�\�B��99��i	�����j�w;�+Aj�4�3]�ݥ�����K��x�j�}��O��/î�ʔϑh]��4���L��"g'��l���kG���7)�[3]q�,R�v���b���?L$(ќ�f@�o���[�ǎ�ܥ[�X�$�����-�=3Uc�$���"�03���7�+UpM�B�3t:Kf�����l��a�ZS`=s:�����n�l��!�Tw�}��gFQ��㋏rd����s+��j}�f�	F=ǜs�آ2�Z�%ʡ�ځ辕�A&'��c��y �q�v�婋�e����~>C�>߅B��N�����YFx��.7Q�t���Ƞ���Rq�9�T�%^ S^y��sr��Cw	���(+���n�E���C�f'�<��%_LD}�������m���Gf����H��t�+�0�LQtAJ}<����e���L���{��N3�SL!�x	4�wR�$�-�\�ܓ�Ʀ�p�S�J)��u(/;�*z��LK�V�a�M���Q�����f�D�UdDbk"�:�)�\���
o�ͦ�貉��(*!�3|�N���|к�*,[1�x?䋪L�>D;ܛ���}Ҥ��z٠Y8�����gq&۶�1"���A1n�j����
���$�+�@�R�aB�K��5ӑ4�<J���/����Nx������Ī)�����<��Nr�KϥT��1�d�iظţa@%���)5
ɡ��+���l��U�_��m+(q�:�K���͖"����̏㹲������lk6)@��6���8
�3f	������v!F�.�
e�A�1@�g�(t�ɴ�`�2�'>8�V2:
��pTX�k�Q����훡�35��w���<�����h����B1�|���O���mD���n�����zL��w��ܖ����^yA�5(�g��ç-F���P���I�����c���C�6�>鑑3�T�}��2�����Jf`�x$Mñ.l&����J`�ū��V?�U-U��;bJ��� ��D,T��N1�� ��@F�ZY��I^"�Ear�]�?�-$`o�J�_�&�I�����R�5��a��#Z�>"ay?0X�8�Y jn5�[9!+���yA��A*�(A�/5r��~�a�O.�t"��kAr�~cLw]x�z���"�Z����Y]8���F�y���Ar�������&ͽ�
�t0�t�����>sU�Fv��
(8�$������/�,����X�k�3;O��%C����/����&F���>����c�D CA�6:a����#RZ�`p��_���q����y#�"A��J8���n�}g1���u�2.ܟ$R,��m`�Ǌ�=�c� ߘ��EL��w�޲�;�]�\F�~X��.� !��=�n��6?[C������PUQ���m������\T){|���r����Ʉ�\4	��:��G%�B������L�vXIٍE� jR;�"_�ϋL-����k�%��G�E��`c*��2S�?sD]��o�ǨV��=�iBקo�i�qA�ǫ���[�/��C��
M�����&��K@�K�vӄEe3g��b���"����=ɟPj�q�t��;�SRZƠ\o���	���捺	xD�Y�?'��ǈ�7e����A���g�b�2T6�����/�)�Y�����g2���U�^�n�������0�f�?�Ld��@a�pnO����*�H�M��������h�C��,�+���'��QA�.:|gO���/E�1�(�i���_�"٬�9.� ����߭�n�=Gq��6�h���U�V�۰c�2��2 ��2G�����7�=�������6�)L߭&{�=04�W��ޜ��02����8� �x-�
���EĎ�/YX����3��w�}.�-Nl���^��O-��F������=29�ʕ��Mϭ-��%?����ы���n`	�1����?�?�H�5���T0f�N�z��{Ñ�X��I�A�e�6ӱh�V�����.�z IIƟR�0��Y�\���}l%��{��L[��"����߬�8�����6�(0'�?Ǆ��K����.����X��2����������2�C�)�:0��a�e��u)���F��ήh�F#B*9��;E���^Q���[�U�;�S�}��(MX� ƽ-R+��J�.;g�/߇��7��V�N��UD����X{�t69��pn��c|R0Rjo#P�O���|g	�M����FϜS"��e�%�3Z�X7���8�����,��ji�r܁��	��Yb��i�j�*����m�#|]!"�Ķn+Z?:�E{���R�����VW<�5Y�J�.������+��?0(e�Zy��_C�2��>{@|�_�y�(t�)%��A���l����q%Xd1N;�<�P��T�'�M��	�l��UM6 �fXc���_���Kkc\�@a�"�0������Cۃ݀-��1�Q���G�X(�]�*��+٦T�s
b۶f�s�mb pG��8��%�R��?�_��1��;�f�������څM�6ޱ�p�a#��5�v��Η�dZ�O$�%{vFu3j�`�b깠0O�`�Ү�:�� ����IK�?7�I�jrHe6ݣu��g�{*�]�b{���H@�,�a&�����U�#k��~Yy0���/]�d���H�������
��5�)�t3����l%�q����f%�c��i�?�u㝦Vid�}X���\P5����gs5Dih9T\���������}s�6[=�	��[�)aO�CJ����3�(�j�6Wty������=.�j����-����ϴ)t��Ir�����qJ�%��s�ud�z���i��G���pmXR�5s��9))TJ�"!.�ܳAF7�.Z��ؓ�4�k.�<?�+3�	��A�p����G��䌯&r��x�U#�]�!��{�(�?[������[�����sq��ܽ0�i��P��<'ȁu���6�u�;-5o�ͷp5��6�-鰮�5�
�4�k�(9|0�Z7�C \�/��Q^d�!�w>���"91�B9�]\T\���n��Fp-�f�(����atc�Վ�a�)����11,h��O���M��&_:�jLs\�j����=�1��OJ���)��y�S���_&S8=$4/���-��Vٲ�_gE�iF��p�d��г1kT����^af75�U������5�@}���_�l�-�iiE��x�=A�<k�>���4�f� �/���`�gd���#�fd�Ď�}��V�)�f� �bzG��(�I��wI�"�=��&�e[��|���-X[m��"�Y�zt��"�������O��5ug��DVh�D�������^'�mVß��$ݹ(�D�SSmx�Ȣ����J�A(""G�yp����"o�yT �$�)�R����2 "����*�r�tW����o�J��#4�9�����g���,�gb�#,�������Z�o�j�n�Q%�q|��}[������u�D���N�᫾�4<q�
 �=���lx[�_��g�Ȓ�������ۂԳ��W�bH�� Ҩ�Cҳ�֏�Ս1�yd��Hv��4���81g�,U�������Ax��V/d�f�=ͦ���J�����%aq��r�2ؕ˒o�x_������ktOc犤��8���K���a9��,�]}ae�q�FA|Yaaq��9�i�3s����ڻF��Hs�vϧ���A��B6��r$eu]�S6a�S�0` ��y�XB���ì���)��t���pO���d�@�N��T��������Zc�)+;��Od�v1O6����J-BHk����'�`*�[K����-T���\�(G�����Z��3˫�˰�Ե��Wf��x���^@���nRt�n��Z�"cnF������ٵ$�i4�.@y�sJv36���38�rWd���'t�]_b���\QY�`m\�
+]l;�j�x�u�ߕ��h�lD�(�z�'���u�j �vZ,��(��@�
�`��S�I����rN����uv�faW��t����zr��T�"0�����a(��iX:`�[$�w~�?Y�e�y�*Pi��H����N��0q@�Q�h�4_���b�熾�[ؚ��8Ej�9�-qh�|���C=��H8}E�&�q`�wk����_@R��l�����]-L�~VtۜR�il)��=Z��n���O�ǅYE��4��h�2,���wl�vHI�W�. Q�j�2ncS�1�� 8�ajx!�� kt.��D�x�3t/�0� �*�6%�>|�R�I6�]͓��§���q����\W�q�ɳ˔&>�3c��IK�ϺH�
}M��s��C��@�z�Bj[[���O� .�);ȣǌ#�jV��{5Sd���Q��r�A�@Fp̹�7�5�M�Ѹ��X6-������^(�f�r��	VԔ�t�@$��&��w-����Ǝ2��'��q@R��y�Z8���{�5�#�R�54�?ec^t�P+ښG�D�'r�o�.6�B��3���ؚ�9vb�{՘Xl��Q�SB�ak���h,��`�I�@�2��1*�F���`(�c��Q\�9 ����=�q��a�-�`�^���V���c£���@��U䩙�����ja��U#�c�j�T��[�j���������/+w����T�mZ[2C����x�P�����@��'D<��m��Y��X\AԱ"t�H}C�x�A��)���(�馂A8��q�~��E!d�Q���L�_��'�]rՙ�Ӆb��MȲh-����p�&�Zۀ!e�ҧ�]��*���).�>p�\k3[�Y��[�{q�v�q�נ���aߪ�'"d��a�W�>����$2.J�3�g��x�~ؗ��@���+�����a^�G� �K�3�_������ iw�0=� )>�q��Y��z^'UfqbǮ�w˸�jq��I�I�[4/�!�!OVvc?H:oPY��R5��T[��`���dᣛ��Gkz�l�M��߀TO��������N�O$f�Ձ
�I�T��IѶ��c�>����x�~�����X��)�� ΋�sPh��1Vm ���"&�3Ϻ��3/�e��ݐEΠ�z*<'��ykY<�h<��T����g��&�җ�j6Y�lѰ�K��|%t,��Al�	���/�⶘��0�3���w>���Ehރs��Qx��`,���3��� �hn�հ�>�ԀIm�VMɐ��J��@�N�K�c{�M���Q â;Mk�J*�?{�������c��2#�6��t# �-��@`^:�	�����U�{�x��D�>����o�i����
i�^�wT�Y�To����Ѳ-��d�� �y�3��%\��<딑z��������o�����Dzϗ|0���/[�9~�j�D�j�.�q]�jz�Q���l&��I.ﳒ�s����l:���'Z$X�D�����7��0�T�QUت	��Uy��� ����u0��39[T"I���s��Ewh��x��;::9d��=P��dM0��k׬!HBag3��:|qZ/?��0���v�3tvD�����+lФe����a�@!fҙg2�������"�us��m��*�
Q'-G�-�6J%Mg:����r:�od[��=>ң�i�#��©qUVq	ެzh�!ټ��i�!��C�Q���ɠ�R�@�G��(���h��my��R���?5MQ��`q���aO��oe��?-[4aT��wF(��r�;J�O�kc��[�R�&1r�}��f�����At�Z������3�cgZ0Ο����$�r��dx�YZ�]���wɲ�Yv��kPb]t��r�{Cqg���D���ie߭��FW�0������<�3xe	��d�.j��F8%x�p��l(�s��v[�D���P�vyu���׾�Gي�0c�}���c~��cS E=�<��l5<�|�͠�T�p�O�Y��X	���?U��/�y{�[��б�D��	��qq��wOK��0_����jq��$j�vdf'#�"�yl�Ob9?����Db��s4���8h�jNa��	:۬A��O��j4�1��D�9�cǿ"���e��E��~�[���
�r0��P�ʦ�}���d�����q��@�pP`�.g����Rwx�I��l���=<J	aaEԚy�Nu�����#;-���Hh��b�2Cw%�/~m�M�R �vٓGn_6k�Y5�Pjjm�2d6Za��	h�W*�̂��������3�V���A��)�免�l����Ya��xGJ��؇]��b���κ�#�3Ws�F�$��b���h����
�+�U�:PѰ�.b#�$Ҥ�������
�l$��Q�0�I�Yz��C�+|,�r����kN[ܡ����0�����҂U-}���jQ
��U�����h����Cm�H�5�&*G��p�����k��g"��_"
�݋�a �+��򪚠���U%�
��a��|Mf�?�Z���	��/?��{Wմ�F낾)���_���Q!p�|�ˊ -��|��R���pϳuH��d��<B����~�_s�k�I����^���ힾ���F?��IF�%�oѱ���]�#k�����P�6�NHr<��_^a!᎙w ����3���(G-b��f�OJ�����C_�Z;K�6p��B:m�)-g����w
��l�D��w��k�]�R̔�ZIU(1#N���q��Ry���w���.��|����i|���B�ʼ(�^��O%Rk}�v��&�ï���j:	��d7Q�X��ZJ���8T0���$r��β����?�=1�MFk�R�wm�*@�W!e�G�9����Q�MF[�{��m�#r�ho��A	>�Tx��-\���lQ?�%��5�W����B\�y9�Y��_��x��8���Wyn�i�)r��D!Ѯܩe�:Q��F<s	I���m;Qnž����w�S�����EN��V��j4p��ޟ(bW;U|��3��Є��rc)�S��x��F��;60L�\Aؘ���%iB�N�3��=�$p*�����!�(��.��5�`�z�L,)v��&�9���ө�3k֜/<�EV"�[N�a�kT@^v`{0lJ�' ������	��=9��z֗�pP�I�Xa$��q� �_��9ī��|ßH��p��V�|�ڢJ������*A����o�ܟK�!i�ϴ� Y����&~�L���F�W>��ܔ�e �R������
���<O��$6�1��������5�D����K��u��<9G��J:���mm^koNpA	�]z�Ɠ�E�2�/�4�$
-��űd�ؕ	g�z�24��������s��Gk��o��!S!��/IPd���x���J!���H�@4�e�hl��z4���j���Ǣ��>5�!}�c�(�@;8'Z{��ΰ(Y�%��� B�[���:�>U����v���B��5,6��Ļ]����k����[B���vm�z�K�����U���W�`|#����1V0�G&�
9��I%��v o�j��l�|�R6j��M8�KX��rڜ�9Z���Bx��%�R+tHs^t�"뉯����ꈖ�md~��үZ@We�o�t�,7�a��XQ(1��,_�	'��V�8*۝�eї�]Ӓ�v��V�)�	EĆ3�4���Ìď|��J�mSi��G��b� ���H�?1�>ĕ��+��K��f�=��Z�6��k�~�5�)�+���g�)0��q��tS�{Mb��,>���H�vmF���D��$*�_[�L�h�Ȉ� �����R���`�X;��s�Y?�4�|�ՖMs�0V�4灗���)�֨/�C}�qE�f����柀+d��޳������1����w��� �@��#�"�0�;�YВ����%�����6Ɵ��Β:vQ(,'�PD���uZ��[�A�(Z��k�i��\$98�H��� e�\B���Q�����"�l���͕��E�IW��!�!Wj=�b����e�c�\eL���i����ٿu"��S� h[��<p��}�K;��#{�g�BKZ�=5y�ҏ���Ɩ���-�<�[	x�Ld�x+�Z��� d�KCW�㵥�DI[�Ο������=^�<v�᧪��S_*tF�� �%�l� ]d������ UÝ�g�w��$�T�*`ɤ`�r�a�&���� ����mH�	���RM��I=���R�UG�sϜ@`���$���4��U��d}Z ���}�j���G�2벤Z��Z"��z����p�{P�u� 7���ЪM*d��M�)��'^$z��f´����G�
�i(/a����̊:/'LRJS8����ߙ�,$ݑ;���OSW~��>V�C��r���6ϳ,&�������H*E��|�G��Q՛�'{$�Rӯ��2��\�5�|j�;��f���͌�����@���Q��w��6�I`+IV%��b�y%2����� LL��:۔�}�x��+��;6������B�sY���|TY�~��S"����I`�ѣ~�o�/ȿ���*pc�G2��:��9/��XZF� ��E���^�	0s0YWD��8��8�G\����6G<1�3V}q���� �Vq�����"tmKC���#yƪ� B�3�Wn�%�<��T��.T��=�Ny1���LW���]�m�E�>Om�����f�Q�߯��w3g"��B6����zG�译݋j�����<p�j$��O��<䡬 ��E�A�J�M��%z�a/#ӏ��)�‫�d�WY��G���)[��K��2'�;�q�=�?� ��J'�O`TeV4��Ƣ=�t��M�^�B��j1�P���,�g�]aґ�o/R~�,DdÌ1�(%��;{�	5؛���L���ML�ӨJ�����f�`2�d0���À���Zƈf۵�K��aoC��(��ܢ\G���0+P�ZHr^�������u�=��U3tc3�}KLע���W��l�Bj���J �\�4h����G��mб�������Q��W��_��k���8����ɐ��3���w,/���!<��*<LH���N�4J�HA�;�є�+�@?���E��/$v�Wk��ڛ��L}ɒ8n�nA��o��u�P&�#��d�P�{�c1x�B�Gt���"*d�u�L���������|r_�����l	��1��Ix|������K�(��鵖���>�u�J�Ov�v��"*و{7��f�5Q7]�#�Ħu��%�
z�̜Ҍ-h�i��sV���ES[��)\�Q��.*�?�w����E�i�"0�a���"�Gk:\����=G��mI���%���4��u�\�nZ��?~��q�7����=p?s����t<�J�����඙��+���SΚ�CE�"�T5xk�d�9L�c"��.R�b<v����;�'Sr�Ƌ��Fr��E\�9`q~GP�M�\�ֻ�f���0��4���x�X<��^������A���N�������u�"}>.�����y��ȼ�$��y��T`�i�c�~~t�7�_���|���Nq�S������0��� �%֭���~�ӹ��e�������S��C+IwF$��`���Ӡ��T�S��|��rX����aJ����h�k�i�)�/���
ނ�m�u0��|BM�^=�$T��&�5�+:��8���୬M=��d�F��A�+Z�׾� �+����!G`�
2����F��z��_ܮ���k�Ғ�F]k���.|�a������� ���bK�!ys�y�f�y@���!�w���Z즽>�J��y��F�3�%
;��Leg7���E��bDoΛd�Z��H?k(�hָ~'Ha$��y;q�P����&�bD��P[�:���FΗ�q*��_4�GW�M�)�����nu���n�.`��{��G~Ƀ>hܿ��q�h&{�	��yqB�0�
F��tt�%p6��{ef�c3��7�u˵��.��J�����(�@�'SQ�y;&���!@�z6(��:��]�8��+zMC<���%�Oz؇�?`�pi�#�w��&֮F�MBT��~̺	�c�q��*�0��Gq:"7C��9�����;��T-�ݰ��3v��DVh@�Y%�!�-���.G��s�r���:�s�e�'8������0:z�o_�~/U��[r�{G{�p!�6�N����TtF�R&V0���%װYq�0���d��W6h��mQ_�ƌ3Vrԃ���}LJ�(�ol��z>��5��P�a%���Bl��f���ba����@ +�{6CNR��qb�/�:O�Er��:��� h���� 7��x�m��věn]���rz�XU��f�5R��k�]R^)��ǻc���n��ܯD��m���ǟQ��1a�K�%j*R:�J��`(�tԋ%c��L�i��5X�͕k��ןfA8~�;*�;����f����t�r�`�㪆�¯,�csL�H}��\��k�ў�2Q���D���e6�'$o����8/�3r���.߷�w��>-qc�+ h&��Tf��d��2�X�E/�֞� �3E�tQ87��b��F���"D���2�!�&7�E���e���@2��!m��q�B1�oh�~�sGj�S@����ɻbo/��`V��C�5P�W1ԛ����a�%mսٻK�?g�u��A7���|"z�_9�q��1ps���Er'�b#�HY@"�z��`�3�t��_�N]go���!�7�hٝ��ܙ���08���XЎ�n��]�q�"�A�a���J��0��� O�7@�l��2s2܃I����XE�h�[۞*�Wob�L�'B[��=>D�~嶃����T6�1�)гGȿ44�d�\�&�d��������n�pw���Z�
��z�v�����Z�VY���������q�� F�]�<���AԀDF��2����?��W�X�Dh;S�.���u�E"ol����k�V������6���C>.�Ǧ���8��������L��5��,���u	���2z��z���c�$����Ձ��
�����T�2�s�ժ�� �z���	N?�?�0����j�� nh�d��<L�f�uVT~%��Ɋ��c�G�xbuX<&���,�x	ǘ"�gC[�����h�
Qn���fp��)Q�uˆ�u����vй�-��Ñ�-��{z��T�S< �d	Zh�2<p:���ID��6��㪖�܄L���G"���Ӄ��7���گ cN(��BJ&�>���J!����Y� �H�KkL����H=S�Z�C�7y��A�ӳ\����-���)�2J��U�'[
"w�E�Ƕ���XE�`���I�GC���-g��J�|#���ƃr��@��䕄��A~��~ ��OYmXli#y�/OcJ�$��)lf�Q&��#ȴb��T6��ͭC9K
_�<�߷]�Y�.��553���%'."K1�r��������	26����2�
�H7�n�B�ހ ��ܠ
#�΃�w~�5_
3j�1l@n�S�����ۓ�����j�z�)��B����"���ftt���{*Hz�[�
��h!��F	�Ll��2L�F9��r�M�3�w3F�<dҮ����'�X�S����N�T�k�;P�]or@ߊ#gauJ��D(���Sw��~K�-��TG���=���#��Qڋ`1d�n'�cA(�xU�y���!e	��m�p�/�	]ُ�aC�Q��=ē5\�2����X�|���i�S��V�����Fs�||�\u%��:y����	�Eꁅ.i���2bo���$㟀*?�$�ԃh�&�I�5�1��]��J���_�����ۺ����+���g�����bq�*Nrc�8�ű�Π��_A��(˩pL�ռ�O�]ۜ�S��K�qS�lJ_T���� �<���l�i�r�ű��z��VeQH��3�vG��iz�[���vt�I�����$�FW@���]�O~GH�?R�_���G���#1��z�M�{��W���z�B�A<U6�	4�����ȰC\h�1�SKYg6&e�ɟ�ag��/7������.Y�����L�e�tv�@{�?c�g)��Y��ZЩ[�RA�@w�w{�<�Z�^i��P��N��M{�w��_�u��7X�EB�s�o�e�vD�� ��X���p#�秚tE^��Y�� ������^�U�x���*s1R��7��e�|�!���~z�ńX�lG ��KV��x�q�9!k[�H�g+��*��3a�{�J�D�vk,����a�pD��Q�j�m�ɪ�n	�-�*�a����������h�	���w&2ZT������<�S�F�� }����$���c��d��32�_��B�q3��_\	<�5�ݷ
�ueW#0��%��ރ���)���e��k_��G�I��
Y����,�Z�m�n���*��0NI���8�l;7D* �7���*v\�J�0G$�w*̘k	�x���^��0ѓ`�P%ry�NW��0ﻭ�}/�d��{\�u=��)�5�l����%�Up��{cW��b<�]UQl왼�U���6+�#�;>?J�ZG��Er��;1��i<�θ-S�k׮g���������8�v֋K�%[�FD�����jr��c���x*]�������� �UxmH ����#$�-��7���ca{����J�Q$	_BN�K�l����a��\`%�$���_bBtS~t:$*�PD$���:L%�z|�,Ď]�)7���������es�{�%��@R���@��@�z���"ۏ}�����s�UU����,Q�W��]����L.v�`:�pt���Sض�i��43
�P~%��5R��&�n�4�\�V���L���q�i��#��Ef8��z?��sZ��Ca�|PFpf|_�-~[��ao28�KX�2Bָiy�N��7�W���q��%&h?�mϒ&@����Ö��Cc|(��I}�4�tv�!#�#����`���JBR��pE�Xo_gkg&~{+��`��*�`��n��1'Bc�yE�J-DY���Y��9�����R�A��i��2�b��Oǯ�RB����F���B�?����"�* �\+��.����N���� �; q /&�sfV\D���r��܊&�z���ӑ���Q����x���؉��̔"��i�G��{a�ƾ3h�?_�J�LEt�0h��ʲ;��Y���"���+X1'��z����C�e�A�����$�_��a��W���O;8s��Y��tC�ٛ9M3�����;�s�,�j2�n�`��?��%�u�FsG�%��<dh���D��
MҖl�׷�x_�R��v@�'��_O�xf�G�Z��n����Wmv�J-"�i6�3���I�ȴ�eN�K�5��&�����*WNk�/�\��;;��%x]ڳ�xn�h b�{��&"���J�P���ɋ��'Ms'��w�U�-с���y�ϴ);�$�n��ڒ�i�@D6�ra�t�:��л�Z�?�����"&�XM���X��\��,���9���pJa+
��*R'F���ͤ�}X�I��6�3�W��x�(|T.��(b>�׷��c�+�g���m�L��0x.�����gl�I�E��/s�0�)�D�K�]D�xԗ�z�@M�_n���
���V�q�՗�z���2n�`DP��2"y��t�`��8�6�ˀ܉��jxb(Π8��b��⎌�ک�
O�"	iT���6���"q����nH:Vz�4a���^�ډ� {��̦^���)t+��,J��!�؜	r�Q9�#'��@�$�[�����<��xfN���n����.p�q�uF*�p��]��(��o�o](�}�����p'�F�T���
�'���J����R:������ZEȀ����$�Q�f䒇��k�Iw����Z�أ9���'7c8VО�$3�c���k��җe^�p�;T�A	z�?0OJ+4cÈCGьה�-�Y���us����w���l�X0ڜZ����1��K�cU����*�0�q���h3Gl��_|a\m�����;�*�*���l�|�;��Ԇ�p����@Z��E^��o� �D��x�E��[�T0��n*�n�37�5������c�F�'����V36'-�U܃+ߦ$�#�� E��,�*�i�����+��+k'���PW���1:�F�<��̛�f��������(��#����t%+���XkU�"r�º��c\+K|O�q%3�PI��.|<Z}u�3�:�s�a�����̯ܘ�cv\:� �H*�����"�M����"�����;2�r/������8X¡����`�RH�ߡ�l���"]�hf<�1�J3�A��ȸ1$�HK�+YBl����]6��sS�=f�}�i�Ʋ����l#��c9��u�D�/LBY�Z9�R3�����(+*�t��8_�=����F�P�5�"~L�L�����P�H�� (���lNbcVhk�Cl��d7�y��-RwL�(+�� �Ա�;���2�ת���A��<���H�E��V���W��̬1=����Q0PK*�!|�u?�@W�����X2�̜wB��a~X�Jq���DK�|��b�PSȻ��"�'?�gn���+l��4�{(�O����9�s�A��:R�^��9�ܽR�U�U��=t����KkT�dSg��h.�{���r��	��Zb����	_�q����/��y��
��Y�rI	�d����PeR2���Uq�F�)[���N2�F��Ά&H+x�J�[�n|�&C��ܒ)@�K^Z��c�Ls>>�]�,���ٱd��h
��޽y�S����9�'ꎔ�%� ���t��T�����L3K���wQ�b=�`:r�C�(~H�;�^�_(c�H�\=����Pxh�v���Ӈ|����F4�)��3�(&X�h_/
�ȃ�W�[�db�`���Z;�q���hL���2C!�	9�1���`��q�I�ӱ}-?u��m�3i'(O]4�{.i?�S��z�o~Ȃ�%fTғ��z�"����5��Y���Uڷ#���E�|ɍI=Q1��[Jm��m���'F 2XoDo�g�_8���.ܐ9�j�g���n����VԯL����D?����,)�oY��EX�Ё�	��n9�
�O(K�*� ZĴ����={�t��,E�I�)�@��e0nˮ�BK����\+c�a�ll�9sO3����a�91l�ɢn7�C��Wa6I&jD�����F�D�R^���H8�=�/���k{wtu�yh&!\@�L��'�hf��)�a���ƅ���1]ã$�ۘI��h�w$
�U�@E���	��ֈ��$:������|�+8n�+��J�!v�N��x7�5�;z"FCtꣶ�~�U#+I����0Ɋ%�n�/Um��XV���Q�'p����rK�s��	N��eËY�cM�wp�.��Pøw��*��;�^����%��6��6�;�DP�aB!I�d�'��H���Vc��]ol����:�,�RT�n�����E暜L�_�r5��Eߏ��D�sG�/a�b�� ��RY�'�ԋT�xW>�5 �r��q"ꏮ��Q�6'p�D{QL�dc�5�ns��N~��Ʒ�б�ۚـ�*k2���G�g�/�ɽ-�16���`���݊2� ⹊��S�� ��	>��m =��0�O�{q���@���u^`��z�J:�頾b��z�>��p3h��x/1�e���f�Ъ���.�yH)ߑʘ~K�� �{�b_G�l�%_w5��vZ���D��?y<2D��md!c����LT���xH�� z}��)[ �Y��*"~�ֽ=}�AȎȩ��M-�>�t�n;�Hg 8�E?�7�b.�X���2(HG5��S�D�K���׋����hqPi�N�|͎�cқX��V|�˥!'�.hǅuc�����D��ϭ�2�DD�gH�9��:A0C"VZ'N�Q�[d��&}��T<Ww������3�M��~�<��c<)�"�N q�|욛'���':f�b���X[�8Z��߬�D�#�N������	�e�̿�
V��@������)ěH��ٓ�FS�����O��f��*�I���N+��/�$?BA��μ���)c��<��1=���kc$��oQ���T�g[,��|j�)T��x<ɑ�6��'!8|6����DS��A�t��{c���4O���J��Cr�
�$���en��}��z�)x(�24���]��i�"�}]���g��=��T�zU�}0����	#�i�;,��lT�O�E�O�~ aq\]��)MƔ�>�N�Y� �H�g)�r�M��k�W�@��rDDÑ^R�oA�kpJ�'©����wo��BL���l*,on�z*4��v9c�l®�X��"�Jx{�ƹ�9�A��<��/ۛ�43X�(f���-L���r�K�;'�%��
�D�& �F�fBr��g4��������nٞ�fƢ���3�W�l�{)���d�F�����Lǝi]�[�<xC>u�~?����m�R��-��$����8��-�E��#1I�Զ�-�QxR�t/��+���u�&����E3$�BEW���,؆�N`���j��?g�:P�m|�����LCŗ"�v� �5w��DM�D�t\���Lk�J��2�AR�k�$��z�?o�p��Ũ~�l�p���|-j��I)R�%���Uw��9�
Q���m/�O�&�����QE��
�V��S����
�{�Y~�]ftʆ������W�o7�CY(j��,0*�o[�����\��<�"��d�eno���W��j���ž���������?�7�+��K��@��V>Xy��Le;=�B�,D�.a�͸ާ�^1�������r"<A����m�6@L~�oK�B���US�$^��aw x�otPp)wu�Ĳ�W�c�TY��=��X�M4u6�5Oј�����RCW+Y���;hLb�{��N�q}�Nz���`�� 58j�k �J���#cѱ�A�Y�
#sv�0��8t4�e�l�Q�L�O��R���v��14wԇތ$���8a�N����OQ2Z}��|%&T� ��v���px���X�i��\4�VR���G���@ܹ���������E��=5U�~i�"�l��>��K˂��](�+K�2iEBS�NL��J��^�Ǒ����(�;�S�S	4ϕ�Rg[);&H���d�:t<M��Q�e����k[e@�dA�� ������a]�!U�-*��=��5D�>9�j� ,~�����'cE����9��q�D�ġ����o�n=�y�(NpY�5�~*�cJ��P�UK�=����%E]������Վĳ���ɘ��}��ar�RZ���mB�?S�1���1
d���CH�U����`����ln�8�Bu��2�Ū��#w�F�#z��A��3Sm������`Nr�v:6�0�6�X1#���À��1ye��I�n��!]dFJ����T��-Er��� ��$�\�I����V䈐�����bV��2�dfl�x��gݑ�V_G,��r�]Q��sz�&'F�|"�f/�/q�F/0<$�;�ot�����Cc�!������1Ƽ7�������������.�(�ƫ��L	�s��T���lfu`"5oX\�Y�S�6�v`E�>��W�߱61~��:ZqE��!��*1��}H&����K��-n�"�91SD,�'�Npߧ�BaK�D7�e+AF�=T횁��kB�m3�+�1��f��
�QPG���7Çg�ȃSñ����+#-�#�C��ߗP�-��=�o�':M�*����Ѡ�};y&��ȅ�<B6!U���吒�7�����@Q�qR<��ޓ'�,�k�C�S�Q��ek�ͮ9<&�hx|t�x��h�nL�XTz�Qj�&zR3tme�-��Q^��K��~�U,_~n���.W��x�	�%׮5���m����P�%����\f9&�Ʋ'vQ�诶n袢/����FK�� u�h��E@��TQƛJ�VF��	�<�䆟��x"��!d�7c*{�	��u���W�S���Ͼ,P}��F�	ޖV�(��IZ�3*�c�=�o�����Y�����M�~BUM���"����հ�Kz����P�)��;V|C��貄��������s�n�U��N�͞�k�I�T��M5�Z��:kV��.ٮ>��q�8Jb�C��4����i��C��n��h�����FW�Eh.�R�k`fC��"C-vfYP���̂���s,��Ƭ{�[5zm��5�����ךT	��!���\����Ǹ�g��Rׄt?��8M�NI�ՙ䔧l��(�=It_����Ǚn{��A�M��I��A��d���H?֌{���\P�����*/T�(����o�~b�9�5&1����jޤV�}���	�-�I�+x��Z\}^�6msf�ܧ���B�c=M���qF�ny�e�6����*�:gn�{���
EKu�
0���T'lO^��\)BUb�S,���*lW��k�L:Qs�M�	����R]��dg0&��f�����t�J{�"͟�yX)@�Y|k��.�D`�g�V�O�M#'��r�)����J��U�u�s/�V��Q��N�]�?�z}����jF;BU͒�)��0g�F�v9FBO���g`���� �����T��Q��#���Tiyh#�6��C�'&~C>	y�ҺFe:�O����eΔw9!��W'Ea)��K;�	\��E�0*�>	�;k�L����#��T<�m�f�a�%�� ��տ���E��a���H���\yX`��Owڼ�қ2��k��]�7~z�G	���3t�la�7y��rD�/r#mkz)*OXl��xy�����%��?��aO�����5�%����U���: 2'���,F�%S��o�gm�9x��]����Q/Y�G�-��Ee����߹s?u0d`���"�v�<$ě�wA�nyM��V�Y�H/�m噛�by��1�1X�c$��uH���;'9,��)�acx�)�*S�K����Y�����o
GS��@抨@5>��9�D�o��������$U|��;�&�WOD8�g��
����7�$�[��J;���p�TGs���`�=���j��IlvᥑG`/ѩ@�G���n?!	Zfڍ��H(��O�Ւ0������W2 ��%���evw����2�����,S����I��[s����C��,���t�g)�j�_��.����U�kK\<�IJJ� îF9zDd\�a��\��{mp�y�:y��3{��p�T����=�wF/�QvV��hyZ��B���ч7Ky�.��m�?�ͱ�S�"��N����M�J|�|��#0�ڂ�H�6�OƁ�<�5-�Hn\�v��j��m��E�'�w	@�	]<�r}&��r���%bl6-��D��?қ���.U,K�:�dn��,���=DF�X���[����$ҥ��������:��p�&2�y�����^]��MsP��4��h ����V`���j�![���d�A�.�JZM&Eǰ~l|	ֲ�Z���`9����]����s;�%������.n�?}8u�<F=-t:��[�آ�L+U��f��@ ԞՙC��_�]�O,���c:������ǉT�D՘3��-6��mj�����rS��Y���:�~�R�Dr���,֧�t���d@p𤾮���F݂�Ώ��R�k�b���=����!��0/��5�n\�c��;���$�Z���1c���_��LK*X�m9#�j��i�����N8{t���9����j�[�n�j
�me����%�x���IInh��=	�sz҉���;��X�ض�[U��R������(�t������s
��:crJ�,K�i"��	�%����@���Wz��j�oo�U�ys���})M%O;�OB 
qh�� �����R�P&�q��+�.w\=���+�7�<�J��׉ԉa�e���sZ�7P���Z[���j�{y\�*�����c��D�)��:����Q�q|��E��.RWsx��婓���e�{慵��G�����,�׼M~�W76�y���fz��3���jb���壞�q�e�u����z�+��2"ł��O:qd���ga=�q�����&:]֞5�����h��t�y�2��Ys����u�5��%ٸ�$�E�4W>��6���Þ(?U]�JA���{� lbpZ.�2W#��R�J]�L��f`NC˱�PEK�[0iQ̍��~�����E�C*�:z����:
g��-Le�O&U�m+���(~z�PX�J��Bq$��>7��f��#?ebS~w�/��f"`L ��sO��(B����6ӟ{��W��}e.؂�w��t���I�'x�ΉF�ץ0��N�@�_���
#L ~����v� �iB4�Xr��f��xQ�w�KhFO �����!Hߓ�n.��?L[E��9/f��3���4g�*�:��`�]�Y�����(0x��'G+�M�B3�b|p�)w�@wp����t�Oj��k��{V�i
�.�wn&N=z.>�����V����vL ���d���]�M��v���&��)%���\#��zW�JR�/�;�eK�y|�&H~A���5����2�mp�}���c�ZW�L��2����-��S'C���z���ݦb�R���� ۹]�ěZ�G0�I�mjd%��-�e�?ٙ�@GQ6&���s�;:�c�����އV}@���I���Qk�z2��R�����Z��~�1|`�hq0�ƚ�ǉ�g����)�(�+iO����WiM�&��YA��9��B|B3s�sh�T�`O�{z{gn�g�h.�65zRy�Pڥ���˔���* ��U[���n`U=��M%e���K����ܚ$7#�\�Ԓԗ���{�qϰ�y�>�-�R�w��Z�}5O�d���}��l�i�e�ha�H^��9_��jsd����{�U4ܱ�6���NO�3	&���^��o��h�ؼл���m/��HWJ�I������L���z����V�g��|�bZo�kOm�*9B�.�쯺�j����-��_WH�} �K���,0_�r�����>	J)0�؏''���M�y�3῭�%9Ui
�ǃ���[<q���8�P븱��+^�6q[:i��?�8��]����k�T^1맲��]s�-�ⱶ�����4N�g=���l�e��k�gg����m��ؓ��Wv2�r_�����m��1kY��ӥ�;��ҕ�/����;`�L�mY�,�5����a�Vo�Q2�> �=J�O��"=�����mc_%8(�PZ��@L��p����KN|b��dW�NW�� {�5��P,:����ˌf�Gkˏ�#��� sS1c֤1�~��*1N.}�T���-��L8.��g@(���"m��6#^(�n ������;Z�����q�o�TJ��)+t@��|��x��8	fH��2�\�/䂎�2�e�ع�D1�9���FzG�N�?��7���,�Sܬ�L���C���?uuR�}��c*KW0�ISM��C3�݉p��V��Z=rA+l�����b����[i�e��fZ��f:r�0l-�;�|���V�f!�xc����y�8G@#ئ.�yGTK�7�6|�����S���92]Ҍ�='�}�cyA��j�)>����$��Yc=����A�sԁU�?w�m���:��L��6Bź�Ov�iȰH+'b]�Q}���
���	�t(o���>k�{��k�Ч(��ڂԃ�h.�IW1N_���*ʕd.�b��j���@��Ry�����H6]����
	�ȭ��,�9FTA|��5?��8��'�����ĭ�˭������{n�墂/�%P@�����2R|�2tX���:���{����
^n�D��l��6%u��S'�!+�HV�yi&��lS�O[�z՗ɧǨ��:h�1��[b�0�/p�3���Fr�UGI�vo��S6�-�X���u�8�����s���,Љ�Q<��	��)8O3Ժ�~9[�p�6�t���|Q��ix Y8Y�!`������?Zu���t6�+�_.{S��'	�u?7u�ED�+r5�N���Uo�*w��~��kOڶ+TD��`�iJ���D��_;�]׀^؏{���%ɔ��H�u#��B���2��!�Wxთ t���� �ngV&d���__&;���Rr��u�IƦ�Z�=���@/{5��ܿh�i�v��wl�������Ub��Uk���BѾ5�Y6{eKuL�J�$���A�9�S����d�hh�2��$*Srj�p�#�6�?ʆp��X1Y�p���#�% ?�~�B9�N���3��~�ܪ��V�L���!<B�!O�i��^��N=kg���rlC7g��oK����fN��f��FX�ӛ��'���+5NŘ\��z��ɰuΞ�܆oh��<�ڙ����Ւ�5����3I�¥7f��%wC�/P݈a��7�����_��O���RdB���)'��_`�Ze1���Lfae��V�����)%3�Z�Gs-ƛIB��B���7��G#p�U�ѻE���Y׋�����dZt�� 'ѝ{x��ܱ�8E�bo��v|�H�X��6�D�0�X8�] /�@.��4�� V]���I����/��������l,���D��*h}�^��n�xI��s/��JȟO�dhص�b-ɨ+�C���Ӡ�����$�q��XH��5�~`��?� �i��rW�;�|�H,V�,U��!ܻ���������.u+a!+h�dߙֹD���p�h���*����\��U��i�է#�=�+�N|$+ �@O���C52�����󑈾¥�k����I���0�XU�A �K'�t��#�?��Q��%��.ihw��z�RUf�E�7��� ,ƿ���.�{i10�'nL���Sԅ������
�F]'�;y`�'[��2*~��`3?����a�h	��wPi[9LE8�i2�,LJ1���B�`�f�n��{S~��1��!�&Щhrd^^HY����ς4�σ��W�h�J.�jk�{�hKj Dŕt�cU�����;
)g��l���}�3:D����Rg�i^���� �L���I�X4���4��|�]�2����k�)U���P���S�/�A�Q����Z���M���S3�;�?I̾����:_�/OI�W����J�R�fL��.����>x�%T~wwOY�u�m#{|m]e��'A����`���xm���~H��̄�
࣒��r�0X�\޶� ��r*����{��T��
�]�*dhP�����j?��Ví5&��.%5e5�����G�Cr��lk-���9�m\�@Qja��R�Sթ��nk�Y���	πD��#���?��V�>Kߺ�u� I�Ć���r��
��3��{�GC�d�EE�YiZc$_�^/��y�3!_x-�x�\��T�LT�L�����S0N������D�䦛-ܐ�Ǳ�0����^?/;58��<��b�F�kݰ��)��~�4�a��}?�	����S��])ތ��$��~r���ce��␬�[�/i!��30a�"`ہςP��z���x>|��;�����,	��S��ͫm��oӹ5)�к�8�aӨ:�O.����WI�����4�6`�xH�ݨ|v=i�$y�ҜW����p��w_�?Go�mBZ�gp��w���?�"&u֤���O�B�c��Rk�H�Z}�Qܐ[ů����ٛ���G@�F�^���I~�ҰZ��j�&�F)�e�u��RYw�G������lK.���ɀ+��ӵ�����mb�rͶB���I�W�Z���@����[��Pg7���2��B�E'0@m�0�,Ѡ0Z��t�.�5x)�R�&\7�@��6ug�^����IS8fb^���QT�t&x;cN��&;���w��DP����Y�K��3`ΐ>�ax�۶1�� .P� g2�"4s�>�X�z�)Og?�r���4�hl��~�P����7Tl\DE��#�-h��������a��e#���]:x,t'W�\��G�%Y��q��z4;�T_$?������
�<x3�yn�j+]�A�b7�F�>p�'`��*���Cto�����4<�jf�O�,Q-���~�=�A�N����@������S�2�tɍ< �ǎ��/��`�����//�~,%��7�%d���J�nP	��P���*�VE����$���}�%����Y���%/-K���/F<�D�h�9`c=_�f:��3�e�}��h6�/������X-������@i�k P��S�g�|!�#4�iaB��C�H�!�M��p���sn
�\f��P�_sﭛ����n#���M&�k�n���/�V|�CZ�{ 1U|^+�=�"z�F�{҉�07�L`zg�Y�o<\&c��ZW�3�8v6]�C��;���~w��<gU�Ʀ�U��RN�B�0�>ސ�$��WX�7�`iT+<i�\��*�c�7p���� 8��[�D��'3��0������:�!���E�����<�Uh�_����P<��ED<�r��ɑƔ�����;��ͩ�J:�V��oj���rN��|#6�:�"����y�ݽ_ί��*�`�dY��Y�>���^��%�-c�ܬ�άF>�D��\t�����˺_�(<�K,�w��g����z��#c�!j��GV�rʴ��@V�+[����w��N�k���~�����}����#|�̷]����:���H�$Ͻ�%<oP��Egq�xJC+�c��I��D��XQP��((�X�jF�봘�/����o�#��P���9��,�Ƥ�	E�]MNʄv��*~Äjk�՜Io�O`�)��!���p�n:���͜�&��JH��s�Vh��bqn����`m��U`;��Y��J�٨	�-���8}�Y�#�[���9P�E��s*H���Ȟʂ��	w[X���R�p�Z��)��$��ȸ5.|쳌�j�}�b)�
7��hF��y�p4V�:�Lq�#
A�4�𠔗Vԟ��D����(�z��� �VJ�����:�5�x�*>!$�@�!�o��ڬ��U��'OBa736�1k��A���T|���+�clUx"j"M�x������ q�����%��@��
������C�a�|�*�+c�m�UT*��K�"��X���8�\���i�F�2W���}{�����B�Y�7m>8�~n|� 7�|Vu;6���=�Ϯ-��櫉��d�55|���g������~z�&>����.œ�&��.�.��A���A�6{P����%���'���>a��s�e3|���?tH�Gf��  ��+�E���@���mEX�����x��P(d��>�W�3m�k�r7��;�6d�C���"⃨�Y�c5W�cp�V��p7EP��^��
ִ���k!A�_W��\чY�?�Ǧ�"�4H�$Z�I��z��M�?Ǟ�iyK�V��2�On$��rUE��3���mЉ��>�w�Or�e_sb �߁�hK0�Q���y2o�K�r,�j+�w2O�|
V��"�Boe46�
Þ0�#Oq�)F:v�S3�d��ȅGWV�Q�,��zK|��7�"�on?{�#���Q���9e��H�l�B�&�+�:ĵf��r_ʷ��j�*9��*psO�k[���V���*���;ݖ����_,N��˯�Z�1~@T�����Ś4��6w��J�s���U��AQZ>q�6���k&��*V*��Ǘ�E�z��*����1m�^sȮ��*�d^]h�qҙ`���#��1l���jH:�rdt'K�qD) �y��A���u�)���J�18���$�Mm(O��<���om=?�%j[t17��1��X�]|�����9��H� h�z��"E0��Ҏdwc�ie���~�7��o��m�Ȁ���h���={�TT�a�lI���,�����E70�nzbI5��Ɗtk%��NX[�Ԕ.������7��CK{�"Z�p��xT҉IT����ô�m,��f�����?7H�F���]A���݄P(�b�Ņ��n$���n���ڸ�o�a�=|�4I��Ԙ,�H��5?�&�?�ʜ���@�_�5�(�\��#dZ	ꨍ�kħ�������1���VK�� ī��jGh��=i޼^���@!A�����N���K����҇�W�aOI��'_�k	�́\�ơ
����$d�vA�U�յ=Di�Q�m
�I��t�D�]�T����݆OJ�!lM�W�t����q�!C��S��I�R��c�$�$�!���u_>,�.�����al5���҉#r=jS�ڨɮ7���b��i*�W�a�`ȣE�����V�v}F"�AF|H��g���m\�@��E��(�I!��mf�h�E�sF�?�y���@�ۗ�o�Hh��Uc�Ih<:%9�Ⱥ颖� ��n v�M���q��}|-��9os���J�l�D����
D�@�fc}أ�8�������?�1US�3S]��	�)	��/���	��A�z�d9RUt��<�<#�QNSF�K?e=�H�w܏W-�W7�^��P�W�rQ��&��n=�ta/�;����U���[��;u��}�5:;�}�q*��|q9 �^>�,�qw��	��
�]r �;Y:Q]��4�>�yA�������y��o1w@��/�	pB�T	���w&�ú�m×�U[C�� �+M��IhzR�4D<hD�ɖ��л| ����XW�����EW{�����kxu�v�XZC���#0Ρ�^�	_�Q3M���	6H�^q�O��(�}���)91�zo_-��љpQ���|��]�/8��Yf�fr�0�,}0�4�:��B9�K�����t��X^��:?9\��c�=�ݮ/��)h)�û�q$�t�*l�~�j������;3lk�w'�֑�����Gj}�F�	���]���2ZuG=C�-�[�+Z/���(����B8U�I�	�n��<n�`\ߕ���]G΁�����(����^4�C����`H�%�播�-%&�F�J��qEKL����>��,�`�┩��.erT)�'�*�&W�&�U�u��2�nNl]^�sa�ϭ�&�^/�&����]�]d�F�cW2� �l>|�d�}.jʰȑ�1+�#kϗ������}��}�[%{B�� ��uMhF�r�����c�d
F���:~�"�R�K�Q! �7�Д}�/:�OM�O��Tө�pz/MT���JÞ���7'q$&���d����cA>K�N�)�lM�Ǽc���pr�s}9�cB�m�48XT�c�F.)^)F�gx	�X��D�E*��+ѭ����b|�Pҭ�Y�b�5x���cf���+n5�sN�B��D�ь�h�)�*�s;�[�&��%�.��qR���٪�i�Eͯ�ԩ�	!+=�Y�+�A��PY��j�:8�]�j=�ƬU�/v5��}��o���d�V���ʈ�Ӎ�6~� ��7}zi�O��k��\��pԍ_r�P����Q.,���%��	��P>�����f�qr"�������$�B]�Q8���l�|�����v��"1���T���:3��ҿ�8>X ���Wc&�(�O�핏	m���T+"l���O�g#�����t���rҽ�m�`�]��i\@���;�lHx���E~U�r.��l�6�k.��j�5%4l+��5e�[�6	8����Ey���f�r��e��r}�8����.��|��h���|Ri4l*��L�<z` V ]��ؗϺ�'l��z�s����_:�A$v�n@X��[��J��ਙá�i�{OՒ�q8>��yqGv�쮭W�v��1z5/��
���o�O"q`�4�f_�'	�70"�#��Zu����GltM@��ՑfTp����;��th!y��<̰v�	��j����r�nVțI��+f;Nt'́����}q
?э�l�j D�H�kp�1�Ί*���t�J�������l�v���a66�7Jc��e,�Ws�]�� ^x�n�%&MΗۿ�Ɣ{��F�g����� S^=�%���<����z�ڧլZ���Y����J��:��J>D�T�2�dq�"i���
�fƴ�O�"'�'�kz=�x�A�2�6;�c�糇�g��ꋢ.3��m� �CG`Ru��/�8N��[�Ư����p���i�nG&��	�:7:#.$9�!Qh}U��ZDKU���<�"��Z����_ N��<����۬�m�-9��
��LV<G@,�W�J�T��ӣ����^"��)g�S���K�1+����E�֐�X;n�Q��푋�E4�y�M�N�=Wʨ��I6���7���CB�l�lBx����dz� �f͙R/ޛY�n3mm6�M��vY	�=��Θ��
*�%���(��v��n�*+��ǩ���q��A�^��iixq��E��7�������+S{�<}��þDo��L=��L�{�ځ��/�SvZ��C��f,AǤ",�n^��F��2$�� ����y�O����}f�^�$@"`���L�&��I�
+��:��A��v��S��6����k%��>���PMѢ2;ٝ�F Iq�P�#�72�^�o��� �a��n�L�C�^�r
�0����g��m���&[ZUH�h�I��?���Fր��^�@�!�:��5�78%j����і;k)�����;�������Z�wm)z!6�8B�U�/�4o��mk4�.c�}�n맼���?�g�c�q;8��)Z})�>;����������Cm��	��T� �Wz�$Q*{�L�0h�\|�;��3�c��^;�]��������\r��ۡu,O�`�R�0��i�0tqIW2��<����ٵ>v.y���%��Ɩd,��Q�G:>���T�x��$'*�+���?@@�����yPqb/���N<]�_{rT����o���p��j�Ok6��q��73��o����OjPۚ��&�����p/����mnW[AmSt�Ǧ "�Л�_��keR���r�ǘ~��׎�ﺱ�٘����`iU7O�6�>�&X���A��{�a���R��ᬰ-	�Nژ��TF�p�5k�1��n-���yɤ�U��9.�!jTװfq���v�U�<|�\�	����<,��$yN!������NT�k3�z�����kX��r��*"~ȡ$%Qk��J�,揯����Ix�+�/����3�� .5��	4-
�:����U� �` �R��5�E�� dYf�3����u�\���;��ө���]G��ͭ5�����*|�m�DC ����&�� O���;Bxޅ�$>L8�]�}�ҁ�[���&�UD�̈�'���)\�XZ1k�@o�b��I��l�7wH�T� �{źoXL&S����J�Yi�</]a(>�~y���������@��[9$�����%(��$%�t��K�=�a����Q�~�E��(�o��t��t����`�����I����!�ãl�����{cG��B�I��K�]�q\������PvT��� Y�%��#dvu�t:�k!�.Y&D݈L���@�����!\9��2\$^�
� �O�0 �x��Nx+�g�A6l;fd��}s���b��J9��:oF)n�0������o���n�lI�e���!��^���4����9[�6�I��G~-,#� �p�_�(<��ܲ�c�S»��2r�Y��?��_�qC�9g�FG��j��"��lZt� ����+wE�N.�:C��
�K@�;F�^;����T�ǭ��H��~���\~�PmZp>�ԁ̸*��C��c.�j\7b�׃�������g�GG�:�g�~�,��8���*��r������/q�Eot����8�n�cI_��>����23
e��iec��R��p�4?5J^��n�B�"�b�蕐H����M~z�"�#aZ�N���^S�RÜ�*���9���"�`b�^gnD���]����M��l���oa�����?�c܄�O� ��&��(!���3&]�������=���`{�S����K����S���T�z4���p��ڿ%��	���T�b��犚�(X��yA���8��`���r��58��KlvZ�4�k��2O��/z�>��!�������n���?��-	J���`��<*`a��VU@e�yK�v{�[)?a#�ݥ���hH.�]z�6��i�M��u�l�2��K	�^��t8s[ �F�P�K��k߀u��$���U��N�s��T�mB���8d��\��ȼ96�+�ꇜz�"��y4�ۮ�-�-������Yz�����<`�90��Dgl���[I��i�F=�[�.}vQz�;��pX+M��A����O��;�vpsDޕ?�PvЂN��tȳ_�25�cp�7�J���_��⨴��!x'�v�#�xO�iF¡Ja�����6��"�w=�9=m�`f;z��l�z�UC�����t}��jC���HN�����I��#��'���p�gb�b0h�ߛ�(�P?���ً�<�n��Z#��
z]C��I���NR�V����T��.x�OV
[0��D��%������0��]���v���n�#��q��A&w�6��d�|�X�n	��~��dBwE�(Yrz�|��/�8�I���p�!
ۡ�n?|F��`���9��]8��Q�r�����:�V˓�����W���#�%Q�{�v<��!aa��sv���1�t��xXku����#�M#��Obz�犝�̫s��M]��rn�F�ꥉ�jd^A��(���>�ry�mϴ6���11�U��p�$?��XT���E
�oN����Du�XM�0�GX�_����/%�ܣ@�\u1��P�v��蓴Q>y�4`��ß����vJ�O�TYu�*U�f�K�B����S��a�k2O��Ka9��ڹr�:E ���9��Ը�^�$��<�w	���(��K�a E���>dv�9���5��(�7o=��c�� Ș$d�{	g�5l��J��f|�=}��)����i���9p�~x�1��+b����h�[D�ĝ������ͪ�S-Ӣy��E9gp��E�Q�Z'e��pY�q��~�T�&X��Y-�Ѩ�r$���UǍ=��=l��i�NA��Ix�(�z�/��L��!�8<�CF�U
��_�O������u �K� Iq��@�e:FQb c��g7�<F�R>%�1V��ʖ��'q>������tZ��MR��hR��r���8Xƃa�(�����j��df���`?� ��ko�ƖYGj˭T��2M*���s< E����$#Y���;��7��B�6�����$=P)\�.�z?^K�����EN��돸��xǭý���zR����d��ٜ����U�o��)j�h�c��X�@�W�65	zH�nz��_C��_R�ޙ���f8R��+(q5�f-�'�:���a]52���H�1����96]�l��am�f���'�4�� �,�0 >�=k�9�Y�@��Gy��?���Z�6e8�\��<�+jz��.�5�UR U$
�V@��i %�dn�G%�|o.���_>jq��!gʯA��k�߻%#,����m;��ҿ�h�XB�ԉj�e���Y�i��LO�5�=le�f�O5��#�爐���H��g~G�i�9�!��ӳw��Em�
@�J-��u쭺7t�j����$xN�a��Պ
��j�A�6)�R����P�(N�`Yg̋�)J���I��/���i�y�|��9�b�Ǥmre�9��}g�b�����5Ց�!��zZe�錇��]fE�t�eS����t͑1٩U�V�E�'�Ǵ��q6׬~�|<��s:��!d�2�~9�yϾ񦼧��|:Eğ��AUrx�3�o��mi_<���}�J6C��}
#�i�<*�����d(NMZ['b6h[O��z�z;����mj�N��e7~�1�v�ls#2d��L����xH?�����q�,�h�'��;�*�	�V�u�
����1cb�u�LgaD�T/����A}�u����s�r9��*�����-�U���X;�����)�@6�ɜ�'��\����x����QTI��,k\��O�g�t�.�K>�f�K�R�"��#��DHy_dq�S+0J��(v���O��^�Xq�~x�v⮻b��SE*�KdZ���C!��!4"�"�jں~��XG�)�g�����
E?2/�)��Ȏ�!�2L
��a}M�����m�.�X��O8t���H��GCKE=���u����kg��z��rkI�"�^R5���&"#{�a����\�;Ԃf35�+�N���x�ɧb���
����BR���#�����nwQ��N<^`7o*�=��1=d�7�J�S8$��\eǉ�	܁=��2/�(����$g�,ՎHJu�ଜt_5A�Qm���f����}DX�%��_��|��OmQ�;J��4�M��Oأ-���l$<�r�Fڻ��m��������r�c��ֺ���m��DxBNuqv�L
��0�+wށ�\+M��k$��`�i��&���5
�Z�5(�f�7K�Q���	$��2�%�a��A�$�A���݌v�8x�Vf�ܴ�j��U��f��q�Tqj�ABu����uf��a�L�� �TFU����wC�(ѣ5�+8CG��0
�|����d�����M��\Ͳ�Ó� �..V�Jw�.�ի�7����<��"�� �2�cy$�P3ҧђ"�ʡ����uZ�������֧_�isI���f��ɲ(��3o�j:\9e
��H�P\7�M�'cV�>t�:����;Ԉv��=�e�Q��X�J�d�{�	��殽�P,�՝$#BC�R�6�����c`��KcZ�o��%��RO�^Z����gD�VWvd�$!�t�[�	ڿ�����w�����hi�����A8���*���J�D�Nʵ,��߃Q!
�rF�2Խ��J�-jt1h׽����5�92-h��i�=�@��QEry��2�_{����ph���⩗5�Y8Jr�����i,b`<����j����6���ؗ�
�M9�0ee�<�0"n��v��=�70��p4��.�c�8��Y��+����o�
9��D9�� CA ȰN�&��q�7��.B���>�0#���^ l|�i{r7,��i7=yk��OT'�6<r5�9�ǲ�5�'��6��ƍ*�e���;�55S^��q:�hQ
|��N�$ȋKUjޢ���_[��W�q�)���g���\�S{+�w��A��aF�>YP56"������!#00dU��.
�5���J�����=>n�6���]oO�&r�҇�;��)]a~�8K��r�F?Pl饨L��� ��M�\g�yF$�L��^_�� ��JI�_S�NTpR�5��1���;����=�=�d'�ԗ���Y�h-rr �����u]6t�J�5q�'�`%DhD1H	n�n��?z�R���|w?�E��)�=������O�QJ�s�6�:�8d�O����x)^!E���iF�|�z?zz� ��o�B��9�?o��C�:B���}������V�
'YB�� 9� Z�ܸ�A.!�s[�'����،*��"1Bb/1��L���5ϔ�%��E���{ݗi�0ګz�]���<�܋X�����n_6$�H������T��]�#5b�lIϚ\��ʉ��̥?�)�4P�?��+"���G~�Ĵ;�ٲQioɸ1��}\Yśߟj����HIW�^���E9G��X~P���Z���ԭ��>�L,WwJ2+�/�FxV��g�M;J������i�th�69x�*G�f����9$�
�wu�����X�s���'-��'����;�v��%�%b�/f˭����;>LW���*>&���eᖮֹ�,��~�_�G��U�1�J[3l7Q�_e�М�CCҐ��O��ꥨ�;�7ǁ|'�	�D6�
!��p�ܻŊ�x'�Gr�d/Xi�B�x���tl��_���R�7ӧA蚇�矁I9�/�+I�.��(�U���$�����EnD�3,����>)e��٨C�6����&8�Nܠ�k1�SC�E�X��z��5�t$�&��Xl��-񕀰v]���dnT� �=�F`�`G�5&X����q9T�1V�g>�������?p9;�&���V^�N��Rfb���Y�#���~�o��+7�_x�o^������ҏ�y�V������v����a�m�;@d�B�nxk*��m�
6�.�����35	YB�G�+�	n�v�۫p;�%5�4G0�KF�x�����3��갽ռ�5!�fMz��Tw!��� ͈��-�%?����e�Q�P�v��RiB=�J=�q�|7����B���>D8y��.�Ե�\�T�f��4��#���%�/FHze��+|+�p�ho��t�i��>���R\Ă<,���U��������Q4j8vE-a��t0�E=�tZP�l�iW��;���w9U��Cd�x�w�? ����Q���������uU�j>a����S��C��5T7�s�&{���D�-]�|]�J��T`?���CW��э�7�����<�s4v�z3������4߽�9H��(˔�:��B�H����U
�Q�ʌ�B)������4��ak&k&�a\\Ew��5^4jb�n�&]J�j ug󞠘a>��7J�Ԉ�>Tdc�c��C��%3�6aI"�����*%�W�*sd�ţ*g�����Ҙ�7�Z�!`V��k�RL'Q�����ۿo~��@�w\7�;�3� M_-�&�1̔R���|�i5�ԓ;*G,�1��5�qPW��Ƒ�]J�?�� ��s���h�wv�8�6 O����eG�:#���I�).�Fn<����a��`�u�1I܋����7��[=dfF^HAN��K��H��8�rF���/{I�� 4s�	0���f�'d�����F�G������w�9���7�u��|�,�s��!O�g�U��j����Sz��vנ����Ӡ��ՓKXQ��ɮ��P�\��^g�̜�"�"C����sY���98���%/?	�ߑ߳��1��&Z�[�LB��L*!hJu*!�P�is+��q��pͺy���
N��2������O4�F&*e�.@����_�w����� �)Y�ȏ�B���WP���p��cL���z
��ŏ��a�b�Q��D�����3!?7��+.Y�I�t��^��?��1`�_��S����T��V#7Ƙ�.ӥ��/$�F��|Z�q�C�3c�y�ۜ���zx��Yh�Z̚����q�8��S[c|0��iG��pqY���E
XUī4|;%_��P#	�A��g����F�!2F<�^���XS�Bhlmh��3B�
�������9σK
���,��(J�]^�Y\+�}��-IoWWH�����j�F��'	M�'�΍>���Dی�gC���X�	H�����_A(����t�%�LD�ު|��aT8Q�f�R�iw��6y�^8��Z]�+Z���*�뻬��t���S�Y_�ʻ���f�XkKY7�ŵ�̏��&���G��m2�=�0��O�aVo��[�>U%TN��뢫!Z[st}�����'�SL5��H��\�����J����hϟq��9±�4�|�Q�_P�jG2�P���`h��]���S��`f&BaQ�3��ѧ�N��MxJ��;�<f�6��˔w�Y|!�+j�Cc�=(`��Y-2�؜^�Q��SO��&�ͮ� &(��	*�K�#f5�^��yU���3�S|��a��)�'6�H��(����5P�H彚���ʕ�,"=�냹�Naތ�������k(���D�[���F�=��N�a=��Jt����J���T��3&t��Bg�K���k�a:DW-�ㄕ��:��IJZ\�E�����!Y���6��1�u7[K�I��l�D�U �����!GP�5cx�R�f����:�:�( !���۴F�����F����l�lر�� U{U~Y�����syq)�8��*�~���/���'���"��1��_�%ǧ����/�	O�����k�4gڽQ�2\Fv:��89��J���f���.U�l2�M�5���_jL���x���S�&��}����e�*ȁ�Ոo\ZwKo`q��ޛ{f4�Zoy�s���Jn�#�/8\�)Rk��n�jɔE��\#�V�k.���'��V9,	%iq���P�����=�`��y��:^�g1Ȯk��zO�p����Zo��&"(呐"�4ɠ]�%���o�B|�zd�~�dw���;?|�Jvs+��R��I���[v�l�M���^��"��k4S�7?�<��Z�{|�w0�!�).�V��$]l�5�FQ7����6Q���l�/��:��J͗0�N�`_wNC��=HW{2ʧ���ࠢ_'�Dw`�N�1g��_O��G����L�[�p�8ܑk,o/UY���g�=�.\�Eq�T�,a�Pɘ�ގU=���n�7�o�X���Q�Z�g�B`�F�K�U�M�C��N����Q�R�"����u,+#%��_��
(󊒆bl��ޟc��X�Ua
&�HT�Ҟ��|8��e�Tep.��6��wT�a�C����8~��^!�:E鍞�9�'s)�J&^�A1w��Г8$+5��7�ص�46�IZ��%s�*������PNn�*e�LpW7b�hu>z8)b&sm"b�㣪`^a��p�<�a�_��x�A��-Ե�5�{��eM^BW�H�J���_��{���K��]�����-"d�^��R/���]�j!C���e��yrHdGӥ҈��5M}�a��ϕ���� P�U��"r5�"����g���P�F�x��%�Ӧ��� ���7�Bo7yD3u�,�|�M����8x�&��'2��>����T��cK��Le�:�S�]�Wyc�S���+���'�gȫ����䶘�!�����a\-O�(�pn�tֿv�H  NL�3 �Ug��.ʇ|/{�)K��ʋ�bf��T��%GV�>B,���#cpj����v��l$�=#9�½л�l���$���T2a0sF:e�(LChO�}�z?8k��@��x��+�L�����C%���t?����:�0|�|"�(X�'ƙ�o�m��qf�
���KH�+T;�.�t"`�f���#"�k���p���x�ZE��ІxG�-��խ���;~�rM�O=o9[@)(��ӓ�S�z�$Bj��H>�$�d!M1@�|l�`"��"�0V$�D�.b��hOp
�<�6���q�\a>U�0���Aw�2�!���G��C��<8���灾���ث��m� `�N>Hd�G0.H���R�T�ϋ�����"@�������q/�pR�>��Za<��8�%�I� ���c	O�5/G��2+7�|�[�ڝ�%�%12ٌ� �c��FE������ܺG�gIL�7*4��-1��zC��?�Hb�i��욄�]T���k�80'٘e�����B%���J����v��Ό|Z�mw1�D��&�3Ir�2��S�x�bx�fqWpKfɞ��zJڻ��I�8����(�����UpH��,|����"�Z)I|01��PPJ��iz�h�7d���P�j5�ǒ������wq=���~Ol�i�g��g��Vt�����y���5v�X+ZK��������'s��/���^ic���27���t3ǚ٩cE��|����7[�i5���:*�Z��N0��MFq�{����I} �F�<[!4ԄO��î�N�7zH�	z��^�R9p1����e󼅽U������ ���/��r��Z����J�9����X4�>(U�$����/�M�M��5B���w��7	���w}��f�L��&�p1�r��Խ� \a��.M��%5:���CdJ7����q��ӁK����48A�V�M�/\a��b����e�+��3� �ę/$i��)��y�=�X��i�8�`)��xp�=�B�N8J���_��A�^���]�ݥhE��ӧ򍺤p2��gaW��ld�ެ�M:e����Ч��\���i.4ɩ~b��e <ϣ^�[�6�l��-+X��t�Kͅp�g�ה�>��X�k�����8��I�-$�Bڛ�~���%��3���-O�#�96&��}��Ƭ�5^�ĺ��;�;̓�������%���%�
Gu�|?|ݓ�+mG ٨�yO!���_����Ϫ��A\##��j}P����_p����Za4}�Z�nZ��^[h:8�Ş�E`�z0�Ź����T�/�1C�������8�J�ҝ0�!�pf-aF�,���q������Z��G~���I��r�ޱ�����t8�o�e�"G�y�˥�dh%޻�ؐ��Z��O%�tDqi�X�Gbr���+V��ii)�5c�!5�m��2X�����JzT_2�V Yd%7��u/���*��� �Ӓ][G/�2�� �Ε*��\��{�"��1�ɰ��H���)�(Edx����<�Ȍ���xx��U��;���Ua�q;m���-M;�G���K�t�5����K�[ڢ�$ݍ��h*!����1�F^�q�֒d���B���)Z�n�X�7�X2_��r���D��F��"o44}�r�F��6�
p�}λ�N'��A��ޓ��������̤���9e0��Z��x���H@�#��2R��|w�揿��/S?1��9�h�x�.wsS��
�ٷ)�	�mț�^s��{Uiӵ�磍V~��i��d�	�����ImY?��lw�\�`>c�Q�ts�y~m�Qԛk�a���*4��b@���	џ\�S�!����h�o��z�N�B�k�yF�PH��x1�m�m��i���[�/Pp ��]SԝL}�j�a�\�(8fB�vo:r�-����L��%�T�JsX��gs*_��Z̞�Q�l�m�"������(��V���;A}m�/���*<ё㬷`��SJ��ֵ���a�Tw���K��#N�Rǣ���GW���M�"0w���2��.vX�gw&�����m.�N�l���Q��3;	[oX!x���r\+�Uq�b����Y���5)Yx>���1������������[�E�M,�0�խ�Yx����HzW��{J��j��-X��g�hX��"�n�,p8����.�"�P���a�?�.s�F�~���}�]���Dk򺢋� ���L�!�DV�<�C��K�zM}ڬ��za\/���[&{�:�{�Z�b��Wf^�l�aͼ��������1�Ӆ�8zZ5b�K���]�/7�:�F�5�w���֙x;AQ��@g-춞kZH/-�^L�(����M���+�U�i�&��ͩ�8�D�ќ�|U[��D,�o{���G%�6��ʔ�����S�(of�|T}��6�F��-V�F�8����k4����N��0. ~�T�ΞP5nCg��j�r}k�=	P�~��36�-�X�Wq�`�`��^��� ����[X�-LS��g�w��h-uѺ�멆��ԡ�V�Xc�e� ����z�k�+bp�G�R��u����6�f8�|�zZ8�E���z��_S��s�`�\~�����f����F(l�y��&:NX��0t����`��2&L�ِs���p�'~]3�z�a��*�jh�8t&z�3�1XP��R�*���x�!_���8= ���:jwH�[�j��Q�a�W5�& ���&W�z��bb�9UO�Jv?�m�D4��7jL�T�}c���y�S�UXυ?#�y�p46"���W�G�x�;s�T���_���4>�!0�D������\/t��uv2������5��k�5�:�WK�<��dD����̤Ÿ�d��	)��/+B�6c��j�e!y���ˆ^�4N�#ބ�yg٦ ˑ�8��N�����ݺNv&/�aܪ3�ߊϙ �ר���-��)9��048����k�r�-��Q{�ƃ	�9[�	*� E1��ڱ01��׳s��3��9ϝot#P��5���b��Y�VH�';�����U�r�t�q���_�/����uZebl�A�C߶������Zyg 1�i�i��A��V�oӨ{7��,�ˬ;+#��k�贴\k���(����.�/h�j(;�#X�I�M!�����ý�4R�5c �3�����Ջnej��+���*%���\�,��æז�BT���/��X&��RhCf��!^���̳���vB����ct�_� Z��x'�c�8Y�Ց.�����<r�+��x�����羡� �p$E�@U!ĺ;E�T|)u���I�/@l����;AZWm�(Z8����PR��zJ;)��V����<Z-�b����3�|ֽ�\u�~�ą�a��>K|�&�@o�O,"������c!��w��rNc�w�:@H��"V1���"y�Ǌμ��3*#��Re�:i,)%z0���8��LrQ4�����_�����i�dI�#�y�Ɓ�����u��gr4�"9=L'��|�A��]hV�V��W
����#KF��Xr%vWfPA��!���J���Y}��T�&4Pݬz�Cn�j��aź9@pf��f�|i�z��)�|/ G�����-�=dQ��(ty��1Ά�"�UE�8S�E��O�Sv�2&Ύ�6�4������p�<�M�c6��ʄ-����%$�)�6��R��+Mx��u~�Yd������Ƀ�O��d��P=39Abq:ۼ�IB*b����J���U
g���dY`�X�j[��ui�*��+ki r���/ڙ�L*�*��/��bL*�^�Jh�2�#���t�S
eli�GkWvY��!vp��b�Qbs���t�1l���]�2�EP�Nfr��L��a�|����1�-�o�����������b�c�6�f̮8�(��9��#��:h	�pV�;��V�����HX�w�3�dV���iKi����p�E���d-�������E&vy��fʛ�2jх���GŗB<0��y�
��^"i��)y��6��Z�V1��|k�����"淂���I����_s���<�g���5$�� o1d��Z>^���"F�+fP�G��t�Z�q�_FP�����i���d+�Ŭ�s˭x��x��Kؖ�O��Y_'ߏ����~J;B� �����8$ע�)��+�Iu>أ�Bɯ����aF[X���\=�'�����*�z������Lw���n�,��.�m�c��8���g����Jn�^p�7ΨG?\�k�%5��_n��*R0)05*��XI`*E�u!���f�8ۊo�i�g���Lm)���Hc×���D��6<� ���d���C�.R�S��em ��?�QyEpbQ���H#}�8�]t�hѩ��~jD�����t6��W3��k݀��z1P8��z��ո0�x}�T!�Q]ˎ� ��L���ʐ����uv/��4h:^��f�`"�Q�*M}A.�h����zʂ�i"���G��X�Ŧm�`�Ci�[➥�kz�f,M��O�<L��`A��Г+uIH�dA�H�?Wc�S�#���T�(�S:�o&�m�=6FC��z����}i�j/��
�A���)�D�L��sS1��2:j(Xob��N�U���fމ#�Y�O$�����3�>՟�p �Cb{�k�U���,�x&��*7g���":*,G�o�f�ڣn����&<�1��NhS����X�C= ��:��l�"�te6{'��pd?�;�q�8�bt���WR��g��~ڃ��tR�,(D:ٶ�~����6��������$-}�W"�˃��!�E�V�)��3�4�U#�����2,�sQ���#�7%�?z7�q�g!!��?��@�ι�1��3�t��&�V"�/l8�~�V`xc^�����w%�c�A�ْ��y�53U��b��~i�	1s
���a�Z��o�<�q��"p��*�b6r�[�L0�����3�g�z_D4��MG�?������xD4GGqh�#1[��e�� \+�B �����{`������؁c۔J�s�@�ў��c��s���	�w���ׯ�Eȥ��/ �L��0"�vc�6�,T,U�b-f����W�V�i0�%�S��˛�������=�.��H1��u%4����t@0�"��f���8Lq+>��V�XU��u�4��kӈ{��� 6��
[ͥ�VE�(5,fwr��>o�W�\\ZW㓊�} �1��\��4z����ĳ���_@}&���.;n�US��1�$�ihLj���_U�_	W��U�N�蝉����EsT`Ӂ����W®��ar���:<�Iڄ��#5�$���D���A�N% lfܱ������L���断�4	�5��sQRk~�۹�%~�<i��Z#���O�z�2s�!>M8|���f�$[���9Fi��Eܼƅ��x���*.��U� �<"�˳�?0-sg���Jif�q0<< x����/')�j����4�����꤈3Pg3
��n��|�E��\r�ھ2�KJ>l��zs������pw��e�76��R���_��`N_���O��
0Ѣ��X���q0-�D��u��q�[{oʢ����X`���;�s��s)��)\oQ���q"�*�_��$�� e� %�`�Y���������"Ӈ5���t�����k�a�z�E�r?ۦ�8~{8 d�bF�R�P��BeƲ(5�����5*�7�oB��ҽI3�N�1܅�T]�섂�����>�Z���|�sBUj=��d�kdźWIf�'�ߘ};A���� �U���3߬�\�#��'^&�t��LV���>����@�l��і�w�@T��N!�E�#s��\u��fP�W��2�O���=x���J��B�個. .��j�[�ji'b�	�_����������m	qו�|N�"����h��UOZ�F٩} q�W/�G"�r,����G^k��0x9��Km"�!�{K�w>�e/=�-�s{�
�S2Um|B
��'7�%������gѾ,̈́<�o׏������p3nc�q�P-�2Z�t�Ng������T|Q}�T������1s���ػ�%ۜ�e��� kt��@�ԱvpcVtdھ���s�R�/�a�u���������]{ߴ
f�����X0�)�+ ���-:U�j��xd#jZ^ϫ�:-޳��t�uc.w��9�'i�59-a�ԪQ�����},�_�Q�-C�j�y	���\/P6cM]��I��{ ��N	��;��(��9GaCZ�mIbXu��I�z�yZ��n���΋}5�)���R	GI��Sv�)�M���}~�	��
���˾Z6�.g�{J���n=�\0x��� ^u�0����QYf�������連��ď���9��t��*$�����\D��A.Ś��\��� ��-�����0���ꎳ��z�-r=����Q:s��K/��z�&�;'����m�<���qBkQ�U
�K�B��n��l�����R��n���c�Y�T��V�T3�˘�s��R�xt�ƴ4�o��`$1or��T�W[�#g	����,m4�YS15G�S���e_�~�L,Ճ�F�F�%���!�|#�qY3.�)�a���F���7k�Mg���7�_KC�@�TugS�����xm����vș���x??8�lKKd,���]^�.*��ɗ� ���*���_��1L�)*��[��JV;64����|��8��rz�s5(`,�|���p"��t[sgC%]�WW�����T �JC0�~�ķ�{���N�*�t�	��8���rC���y��Y2��ʖ�5��*����ݱ�-���v�r$�dp���vD�V�n����7'��&�Q�ؙ�,2ƹgh�iF�	�&��O,'V$�[���UP!��6�/z-_. ��X����kjnQA����UGX��=�o�^�-����s3�	�4@6���g�gR"����H�	��W���]R,ȣ'��+a��f�Uט�)%�(7�Ad�p��!5��\D�� Y#�f�}�=J�Ș�8b�+a\T_��\O�_���'����E$܀�~m�s�i���="���׌|�3��,�A��I��t8�n�^U���b= ��ļ9�Et�8)�,%_��H�ߺy;%~�n&����-o��V����d���A����i��i�9A&�s<������HeoAQ	�DC-j�j�d?�@���̤�כcTΆ�$eђ��6n��m������q�i������5�:�t9�x�K����e*D� �"Y�]HGc�n� t����x�w����m�d�rY[�����1�푬���T�K,h܈�8G�!W�`�32� �f���VҲ�ן��Y�Fv�vz
�,*tI*E`2�[u��{Z���?g���n���d��]Sj09�\�L�^��i2�o �ٝ���D���;�0Gk&eZ^H 47^����~��}���f��_�w���@yW�C�!�mv�������L��[L{���:dǃ	��Y��5���xwH��P�A6������Ïj�,r�u�]�Z�1c�2����[W��O5���{<br*���<��p蒘V:�s�.���鍳�=GX���Շ ���9��K���'&4Ϸ	LŮ���~��^L�b*�])����$|M�w6s������6
�a<?���˒6')�JV�*¤�5���p^s�][����Y�I��|.��m��ds�RTW�P�nQ���oUA��vn�X�KJI�14�X�|�FpI~��DVC@������^�-�6�z��tZ)��;T{t�Eo"H��)��6��a*h��]�C��%�d[�?��a�A��FF�`���
'*]
u�y�bC+���y��
߅S&'�.r:��.�ެ-s��^�EB������o�����7�hJ��402,�l=k$�b*��b�� ��S20Ys�4�f����ͭ3���L�S�[�o��Z�Um�TIT�60 ��x�,����m�?�Q�ǒɼ���UL�����V�f�p$�Ԕ�>�+̗L��Q6��t��a���ʱ�gF�5�O�W�ܕ&�����US��j�?�1����a�V��6!D�R�i(���zB)�q�~��\��5qq�(�\��<�� ��#�jتRX��#��]ߴ����x����!HG
�?���G�?�f&�Xx�W�+���y��fcĠ�$GB9|e�^�ނ��
���k�/@�\r����*\�I�z��<&��Bdy(�;�����!Z���I��ƍҪ'�`~ge ɕ�S<F��˞���7'�<6ZX)0@�y�r�X�by&�؈M��wW�A�!zb]��4��j�x�V��"l���s�������vr�֐?v{lo��P*�I�<�s��kt쭐�	�(&�H�_�Z9�,]��3�Π:�gc*��0 "Z;[��l�7rN�B$�H����<��"3b�I��MX�|����G��9�y�Cflߓl�rNy��P��炲��<}�;�ۡa�v,�[�>�`���9n;����R�Hl����+��6r#�I�c�]��t^H��=��hգ��J�4/z9��˪ip\�۵/[w�������߼M�IP�y3�0�sBѤ+�����N �K����5u�Ҍ�$4�<��E���\� �����obg��y^�Wa_���r�Okg�_�����-_��l�/��M�	�൐9�6!�%T�2A���JPE�(��� V��	E57<�ggu��|ݙ�z3,�	,���\ dA�@����+u�OU4����ә2Q��b��{���.6���F��0�O����H�2Z���d�R&�S:��dK�0�['[�;!����`�q�#���q�!����jY��	J��uQ#eǌ�+��Ă1\̲�^K�x�ۃb�j�m�A;4e��,z��g������Ո��a�⨕�l�G�Sҕ޾�Ns�>,E�
ݟ��:���~����d��G�un��[4U\��v�	�	���v�v�K1#� ���Hd��X�?���Å�wnv`tg5@RY��j���;bfڶ�)>�H:�kaiݚ�`n~7k?X�P-��rr����#�1�[Y;�۪�{�jM�[���AG��J�g�Yu���	�W���BQ@p�"�1�5��� �t���W��wZ�|.�_�t�V�c3-g��\齤���_��3�&�2NCB���)����]�)��U�B�`�˖�\��O�<���[b�^v� `r����a��,{I�C�Y��#�r�H$G��;��c��5[ڥp�!�~�%V'f�n���O�iw���	d����4�̆��X@���ۢɺ�A?�r6�ɇ��pJH���HA�k\4�ؙ�I�����%Ku�:��⿐`����y]5�c�W�$����@/=���n������<?a�>2y}�Y3���7����Ax$��.���Y�y0�)�u��7)z< Ē�^yj̓��{R,�[�I>�[U����Ăd�������1���|��7u^F�H�mUX�%b�M?�d+���
�0?4k��Q'%�ͺ�j=w��7�$��~=2��^2�/�Y���]��Z�N�~����>�J�c!!��ee�'�cH���W�䧙hq�SJ�
��ɟN���*4u�bml��V*'����V�k�8�lnZu?S"_ui<��
mؚ�*��S��P�(�|�u '^i�|MH���Z� �[݂�X ͽr��t�rڗ>�%��[��=���o�+ ��[�7��0���A<8�C���U/����b��;��Z	�;�c�#a�w��.��������m7�"�B��_~��}<��5�:������}������tLK֌��˔)5�#��Ͼ�A�KR����WؠElY�u�d�x��3���8�KDMe���,�z�"��~u6�2r����v�䃚}8	x�U)�G���߱X�܈����M�H!~�Z���:�~��7v7[Z�d.z-��S��)������jm�RK�qd��0����13�~^�k���~�C���hk�I���@@�M��\�Y�`�d.||��@޴&P�stMm�t�9�@���脐C�ѥ���΁�������,�{��D�I�y]�7c��It�ӃxDI��]x�Q�1�qI;*�`��JO/$�5O�s�?��_	�04���-J�8vaV���I >f6�M�A^on�/s��k�GS���Ѷ16x�;���5�Za�[h�n>�O����/�m@C��Z��2	粏8�`20tu}lr��¨k2I'h,���{�u��g�����B���KFT��ym����������ƾ�*�{���-��־�m�TdOK�D ���]�~y�M�o�`���ĬDS���mOy��з��SU=ՏgtW�^9�ߛN�K׆��v��w/d����$���4HȜ���=箼��1+��' ��,K7�H�5�K�ic1Δz^}:߭�"a���W �Cr_��M�k�W��������a�\����6ˬ�Hř����`�����L�)�W5�(��̞�7��n������F0���MR�B����S�S� AB��V-.A:��\9�&DO�^�x_vE��i*8$���]H�U��
⹉v��D�
�HJ��a�@�dU���,h�xOc��|t㙐țk>χ��W: I4b �A�'K������'��<FP��[�i�`�[���)�q��B��q$eo��?GN�FSx��X�uץ�_�Z�:|U�Pͩ�E�C�Z�,H��df�z�3�e-7�^���6�M��n5�W�H�~�M
Yd3�lu�����:#bZp��%�������yHhf[����0�����l�rir{�d����B�њ^����m�o�R�)N3$�>�n�\㧆xl���*nw7�,@��t^�G{����m�̳I�b�|�L��Oj|3�������	y�����19������[D<��WF�)
H�.���f7��e�U�E��X�n��C�O���ޫ}|׻䎛���,� �7�����˼���{:Q4�d�tՋ_���땙9�����*I���B + Ɔ2���9_;����c�v/�'��[}�ˍR�R���TyzS�k�>	ַ-���ZG����5�6�r�m��P��7Q�o�{)�����<�N�Β0퓻k�p�l�Sp����Q��U~`�F��|������V�(v�Q�&ǳ�v�-�e�å��)c�?�*"��)|��i���)`0Xvh����ѭꄹE��c�W�����p�z��ɬ@n�Ԗ��6m�,E���[��, Q��)��e���.�h��*c�!f��4��36�D�˦0�D
�9�b7"fP	�c?=����3IM�����^��1�����	�?d�JwP�b�,��"��9��'��<;��
������ X�Ɛ�q�|��9�!�"���"���nCۡ|���7*ZZve��WV����s�bx>�b�����!F<������qtvO��n�^�A+zZ�b�A����I��� ���m�7\XH�#���Q�̆��0ݦI�;� �j�*��S�[R¡ᔒ|���
�}�f�RhY�%�[r�9�+V'+ Q�5�eҮ����&����gn�}'n�_Ŏ���1## }�n)ت�)g�0?ΌEH%�cJE�p�n8H����)n����t�`��X�,��oZ������#q����_��o$p�N\��ShIխ~tv�7?��!�~���n!������~cc�֭�EX��]�d��� g��{��E��ݩ��r�F#�;c���=�x�� yM�0\C���%4�	-���o!-har]�FJNs���.�+J�� �|���(����W������`�~7�hD+ �@��N:34!g�\f@�?�h�a1��Vo��V��+��0����*&-99���C�n~]���l�?e�H\::���#o)u&�0)��r.o�E�_2�� �=?gw��R�,�[N�t*r:�U(Tϧ�����[6�_���! ]Z�]��=ʽ3z9=����x�"q��1�f��]k��	�E&|(��k	%���`���|_�r�D�>�����Q Xc����>�SX�ﴍ����~�J~�;�q����	��|D�e �")cF���bٮ��p"��� 5§D,k�U��*��)k�������!�=˴�*0�E�7a���>�S�k�T��D�6��=�\�v��P229�  ==	抩�yۤ����z�E��� ]�L�EMQvAFyo
wx{��L�3��i�u�vB����ڛ}�U��	��y}�Ɣ�b80T�l��@���V���ؿ���k<����փ'5��o?���(� I�
 Z&�d�C�Н�B��*u]�+ħi��>�g��kzH?��d�%�+E52Fn�!��)9y2�?�P��t���O�Wշْ�cQ-�e����|zq�0:4'��|���v�}�3]�>;|�ub�d�������&����{��7����XPH&To6�<�J�O��M���jGj�iNq��2�n��RZ��o���)J�=�<]�_��x� e?bhi�(*�]5c��wq{�L�h�c�"^��:��`E��mp���60�LX��ΰ/�J��K��B,����U���K���^�uk�HI����#v���]����z_p�YZ���+ڰ{B��E�` ����*����	-{P��a^?�ޏ�>MB����%v�o`�����t��lN?���f`&���u{$Ñ��n�`P�n��;����̻�'�u[Xݪe�(�`���T����m|o���yE��HWVR㍒
Zd}�!�Q�zCg�l#鈔�[G~3�vW�SE��s�2/�F�=w�к�m�|�T�;̏󅍻y�����tn&"v����d<{ �O�<��|�G��HH�3����	_\�*�i� �6����Z�m�E�J�d	{U4��1�K�+��Ƽ�����Kp�h<�Tm�����:J���� +q6��E�U��p�	�r4:��O:����k�m8Q!ɺz���t������Vbg�U[��m;���(R�T� ��+�V�
������w������Wb��H���J�x���p������h�@����1�mv��SMo�5�#_�01�;�w�m�j���c�QK��`�G:�/l�~�3M�#��@���$���}S�F��Dw�C���\�X����)fw$�i�k-+��j^8��Ӌ�r.�w=*��1�6V�Wq���Y�΢b�>��y�o0w����)n�c�;\պ�(���w:2������)^NUɷ�b���d��p�y�i� ��~?u�?�ޅ ��#���{
"i�ەr����|�/ǚ��>�vw\��?Ko�[�j��ӛ���Z�&!Q��k�L�S����Q�"�1�r_����L1md;VW�N�X!R�Cn�j2g}ӻ��3d7�?�'$d��<�'$'۷�Uj<�9)��p��@h���|-�@3�����l2R.��Y�[@�����_��]�L����ש֦�A�����IO� �j�12���_��!�S�n����(�����f{��ㄎX3��S��YJ� "��LeK�ȼ�
� S Um��⒲�,����tQ��:=��?;zjI�=M�H�OT�'@�uݡe�Ts����і�A;�Z�7�46��FX�����ۘ^oH΋����\��RȻ�6�}��G/��-bh�XTv��v��ƾBQ��sWx����k8ᕨR
�x\����!V��i��	ĘRXD���D2�2��t9���i�~b���g<���q�G�$!5`�h��Xx3�jN[�cU�Ni�Bnf�NG�oÐ����S����w+�.jI��V;��^�4��bA<b>���p�H��F�-�����\�KKx`��p^�DX"3KI�"p��h���T�m<�2�Nc�T��;�?)�g�E�I�b�����4 �G%���*�-L��eݘ{����	�R�M����I�T�s{YVpU�SMǅ�7��P�)�b�+4t���)���H�a6_E���'�Wz��^���벳��muY�Î/��&_nM���q�X����`��-���$����kD���W�~� �V�;�^X�=�b����O�-,��@�~�K���,�Z���%��:1ֲ/�M���D�P���x�pC���r�=͒H���e�j�����(Zd�Q�J�Ф=��P�+5�Tط�b����w}���A�|T:����\��=�aY�M�9�{}��M� ���Ԙ�{va�"�}l��Dе��0��L��_��5����D������D�<�; �`Jk\q�3iS�#V2~�M#Zȗ�-��Ő�EHV��(6�R������M�,�t<5��H�33� q����BU�&�*��1����`��h��9�W���Nd�mx������DgU�:I���)�9��H��L5zʘoB�E��'O��D��� ��s� (+�0��D��K(�y 8e�%��J��^ ������+l�aL""'�2���zU�QlD�X�`ע-�^vǘ#�����<�u�V�Թ�qo�M��%�mt��{}ָc!%�P�z�ϕ��]@E�4�>�8����*�O�Q����%]"�����|��%XK�|��@�]P��)}�Ā�js�1�rOQ������h;7z��`����{du���N����1���J�%��a�4/F�֯��)�C:�7g�r�R<wʬ���²��6$���6�Ӫlɠw�P��-���E}�M���g�$Z-L�	�B�g��G�K-����*8����[�����؁��{{���(��ěi����H�CTG��MH�F	e���W�b<��~�CgЍ��Щ
�w�Ǵq)5�a�	 :r��RT�������# �@Oi��w�|�!ݸ�]x~�S�ћ�� `*�Ӌ �Y������ Y�������������U��{���7��[[jxX��~��T�Qh�E�k[s$>�ɨQ-	S����/��b%���5��Q݈��j�i39�xG���=���I�L�U~vCd���ʠG~�] �����?��ʹ%B��@1�H�:�F���[
���/��*ס�R-i��l��9ój���X���#�68|��:�����Y�t�]���Fƛ���q'�=Ɵ�j��.�}�o=�?Q�,���I��M�*�e�U[��j��e��91|��HT6,�(�dq�^'J����R��p��2�ֺD�0�  9�v���a�'�����5�CuT�TCy4vyR���6�|ڌg]4����i�)'���d~�24�)#�,r��� +�²�;��0i�$-�������L�5���ңQ8�d���5�"��L8��%�f�3�Z�3J�����fz7�kR��J��j��@*`0u|�o���'��;�h0�Za�(�	߈�9�c��I}`� �}e�N	�
�
OH���5uS�I;�� �D.����|?I�Rf;��B������M����"�h�[�(4��Lm*���L�Q2Q�)K��sb���q_j���L�%֔�ifh0 �F?\�:����H�e7����G��"���2.��PX׺�4�m	����s����P������i����X��	K(ۛ�l���9?���-����P��}��6��Rϣ>@VѕPu�-%"�y�D.�f��Kki�%Ծ'�R;CQ�fÉ�Xa�o{LG�~`
D����� �[P�8��h/Ż�P����g�@UUH�9��?�/�f�°e���:���&��=�ٝ]My����<�[Ȕ���,��L����@ W����a����Ͼ\?}`ޤNj����DBm,Z��y����۝;�<|��5x�r�C��my�G���#�I�ٖ3���q���f�( zS�ˀ����T��<,����Tq�˘��6�tO1$�ܑMp�(5�vm��)�{Q���uG_���^�<�R�����+x�I<��8r�Q�],�',�	B���:0Z������z:
�})�����$�V��^Ն�������߆�Q��*����Ҋh=��q��-��	�-R�����2Z�	H?0�#���0/1�\�`|�����1}ԡ�hT��۫�z�Vy���[
I)dA��?����d��3W�mo�Ἤ�?ǫu��%��໠���w��.KhFCW���i;�$>:�G�L?�=XZChζf1��R�^���ɍ_�C3�t]�ʆ���7�Q�	o`w���@�xE-��L}��*�Ygo���~��A���y�� ����twP��^�(p �.�i�����e� ����$K8��4�Q��<����KC�!Cs��O����߀K�a��R9����!�š��VS:2�"�Vl��7ϐ�(T��dp��y'Mc\�������:�KbhP�K�_���;���8�bx(���ȳ;�Y��Ȯ^m��tjݜY1UҾ8Pl��75��2�3��H8 ?�=mʍ�G=���nc,���;
߬��G�˝��J�o��飱�������M�qv�_�����"D��
�x�rk ���D%`��\@�/����<��z1ͯ�^�8f�%`�"� ��H�]w�O��s|���:��W~)��}&�5���]nQAsп�n�"�1ܿ�����!3�ᖬ���I�7y�%cݪ��5c\4v�@�}�3�D���Ω���S��*ȷ���ӀO���GK;�i:��Td#��EV���}��;�UF�ѕ����8�*�pq
�н�"�y�Tw��!���ݚ��Ւ7����/4����]�<�ÒX����0�:��m��Opn���&��5����+��J�]��Ȇ����^YIC��k��Hީ�=�%�k��"��Y��۳�fGF_�b���'_q�����R��A%3�叹�q9]���f�v[�&�9����5)Z���Q�s�缥-|.cDw�\%���w� �w�ʍF��u�}�mǣ5�W˯��,�x����@w(Q��Ч�U�^�.�����?UR�-�9�\��xb!�%�5� {�sip	����=������J�>Ϭ�X�g��!�����X��2�M|�k@���V���MBܺ����{9��=��A�������Ъ<o��!�q�]j�P:���l�:̳ �71���7:$��'#t�	�3^��փCSh�J��C��i�F��`p,���~{(�~�W�O`�>l�}��E�P~QJLW��Z2��'k�IG�޵kym"6�JUκ�h�Nh=^��s�Bk#�^����Rŵ�hQ�[�h���ܻtQT҂�]�1k�^;3H�@�����T����RĝEi)�;��@|v�qyz�9m��뭽���=]Z�c>�������6s+X��a�/��A}��Iɑ��۰g���duuW�S,,\��-�]�s/pL����|r���*��A⭜6	�����-��Ώ����sOi?7P���8�J&C��e�ź����j��-OcUh��
U�3���9���^�p�/�/3�BX��f[}��&W���ϨĬQ�#�h�`����\���/�7qCE���m]��[�%g�	�1��6b��Y����>Y�^sR #!&�w��11����d�;�Χl��ArE�=�{�!��˭�j��_T���3i����)� cv�X�+���?.R����o�FL�_��jM1{#��!d,2Cb��iO�c(u*K��3�-�ϊ
��tǌ��G4�M��2�ļ�����OåL��`0һ��o`����jT-y�p���*2س�(����{������1�3�ui����j֢�Q3<d/;D�ӝ���\��� V�\��j�	�������W��i� (���r�em��ܰr��ݎG�$#����_���K^�(��P~��?\�ױ	o���&�]�5�ƞ:, �ܠ�z}v���a[�* @��Q-(���ʃ�����1Q!��͛<b�<��2y�����V�p�l�x�O7�2�L��V��VL�4KK��XN�W��P9W��M�Ρ��v1K����Y��ၔQR�8�n���
Q,*ȝ���`(b�fRzN�����V�Pdb<~�h%ѿ5G��<O� �� �xF�Eɂ��Ɨ�BM~Y�����0�|bxŏ���M�dW�K+)&�(��~Н!�����"�oF����m2�&�Y�A�Rl�����)�+K�U�	.c�w�K:�z8��<¼5Ų-=g�=��0��� �� ���?��^�Z�����Ak׳��F�L�k�����Qx��#уbAZ-zwШC�_�5�8�Q.ⴙ�ꄽ�7��::{i���菷�9m��� g%��AgS�ju��ȳZ��b5����Ӭ$#R�H���v�d8zp�3����
�13Chg�M�w�u������
��8>P�m���Y��}�{:���ڰ�og���XXY�>���$�~�e���=��^B�����N�D߂��e�+p��e�Zf���k������"a��4/Y�����J���zi�u*[i��H�{�����'�ZŖ(k���T~<d�f���$iX:0=�`��+��僉ۇ\)$��x,b�K��y�������7K͊aIs�C��� �Q�*�W�8��w��p�8�O@^�"�Hp�h@Y�ȗ���P������ܰǹ�x��Q>���;����Rļ�WD��]�qcƪ���N�*Y����<�p���:th���"^��T�Ȥ�ۻ�
� O#��s���r,�9�Fk��yӶG&r*��.���o�B��zy�~���$eO��i�n�O\��� ��J����;O��c�(;��K���򵙡w�\���ͷS����vT���'��{m	T���Q�mkct�\�a��	�ۀ!_��d�*�M֝n�uG�5���~����-'���P�t�̻k	�ʷ@BqnٯMh�`�,�
�ٛO���J�?�'�R(#���t�H�����Ш��mu����s��U�/Iq�G�$�e�H@��b,�&�k(x�>���#�f�ov���0���g�=��lOVsWPD���%�qz,ޤi�`�Ё��ٽ�1�d?h]+x���@�����+���&~�K��hc��C|�QЯ$���~�v_�K��5��'d!�	p6��J�����D|�a���ō�f��P�:|��7j<�����6�+�RB�kZ����+��nh6�vF��#}�vț|1m,Ņ�3W���'x�c<��˥�#G�&�4�V1	�>�ļ�
���T��ùtN{HȮ=��YT�a���"���G�O�"LɃ�����R�n�����F���&�G�Z���m�;9��\�)0"���[3u��P�ŀ�ˠ��4�l�����K���h֠ps�D�V���؃�4yFg�{�c�X���!:|$��q+O�5���[����6QcJ]�ƠL�_)������(`%��FW�Md|���(���/���9����۝&'�yEӗ�J�N�����q&88��[vq1�3�$#�cS��݈��~�؞��zZ^�xo����9-F5OQ��܁h��r"\ɓ� ��Ҹu�M����m�#ž���f��r��������_Ŭ�xu�$3J��!��~�����,�r��%�����>k�<���8	�	"ZH��ޮ��%���a����*%ȈHp�_����i!�����x�M��:E�/K��c|^)H��Y�ts��L���M��ò������B�����?�1��ɋ���_d�k���re����L1Q��[������I� �Ya[�x����?�g�GK�:>�H�c9�s��a�?ӇDL��C��1r�x��g$�S�����A7��Ą����͹$���1�F�"d �Ǘ����(a�td�(���T��e��ſ�^�}��&��<��_}��:%�����C�D�(�f�Y���j#c ��
��\/�ܒ��6��	^�ϤĠ�*Av�	��H�p�k}�Ĩ2j�x6m6h��Tĩ�H��i:��޵�"$����զݟ�*�O���F�;�9n�%K
�ȸɥMl�q��Q"���ƕ#�?�ph�v-anVP�&H���F���){��e�e�'1͢��u�ʷ9U�^��t�� y!���@>�����p�f��H���ר>)�L�=蔇���Y"Y�A��(!#�b�.U��e���R��yHio�:�����N%���W"Rf��N���	��mv.�W�z��i�EB��ymN���3&�T#�̐	�D_b}���GP��ha�)�k��m���6.2��r�"!q�z�Vo%	?��^2e�AHkBO(|sD��)|��X�Fqٟ%d�[C �2�v�S�����zv�AV�+���v�:Ž��]�(����\���=����V��������58?qAц@�w�u�+�J�x.�`vB�O?X]�Ǹ�Kqh�]���qσ�'v�&Oax8d��#��T�����_y3y�~�C�a�h��F󞬃:�k���+���lB�����|Erڮ�5�΄cǳd��AR�zpA��	&�
�?��k��	��jvT���
^����p��>)V:����k6r16�Zcv@����z�"�֬��HS�K]�m�I#���0�w���)�� �����3�A�=i����G��`X\U�:,��Y��H^�l#=`��B��i~QE��$#�*�)]�*�~�b�l@�e��_[�	����j	~>(�<{Y�߻ZH!�V�vB[,���Q���n��� ��'4"]ؑ=�x#f7qt���y!�I�Jje�R����9�*۞8a�s�]��,�/��ħAQ�v��@��"���6�E�4=����u�IBƯ�ڳ#y9 �F����	�K}���G���"��4V��z��|`�ЀN�;��dN<�M��O,H���������zR�8f�YFu�kF^�>G�v�?R)K2�,��׿��@Q�e`D��`�saK�8�/�^���sr�{𲤯Z�X�������rn��h�q�n(�=��9ܥ��P�� ��'L��(e�|^K�!$7��KF���只�����B$�_;�&�'[��7��a�U���0�9[w�T"�X��\�ę����X�j�X�& 7@������k �hn��H�W;����گ����guH��PAv�<Q5 !�
��V��� c.5հG�s#�D�a�PD�̉�{�;���a��`��^��[b�&��'�q�� ���l��-Ӑ)&�T���պ�Wӊ$��G�Yh"ǳ�R��{�Q�k*�/H�8U�mo�fu9VeZ"�,�=�|�ڪ1���/�X��Àz���ς'$l��Y�+C�f������p�s@?���?Ǎ��6 X>Rq���q���έ9��7�J�g����]����d�Պ���"r���g��H�"��y*�2���!%�X4=��m��o�T~�Єs��.9TB���>����6Z<I�5� �������]������6�S�^8��Hzu3�i�X�<O��_
�4J��k�X�T�%d;��m;K��*���a�Vf��]�z �7�i�� ��g6���7�fx"������.\{�v��|S~��py��
�/�qopd"�m\M��d�C4�9cmJ��w"zt	�V6S�+~6iԚ�(��e��4����>�Ve�A��w��M�Quw�8T�	>�`6L3cu��#I5�K(q��)t��(�2����ݼt���'Y���t�F�b[vf�f����缳ѣy,0���b��%�X7�̤Y��x������ ö{ս�C���